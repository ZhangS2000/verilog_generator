module sn(
        input clk,
        output reg [5:0] led
);
`define INH(place) ((place) == 0 ? 4095 : 0)
reg [11:0] p0=0,p1=1,p2=1,p3=1,p4=1,p5=1,p6=1,p7=1,p8=2,p9=8,p10=0,p11=5,p12=9,p13=0,p14=0,p15=10,p16=8,p17=0,p18=0,p19=1,p20=1,p21=1,p22=1,p23=1,p24=1,p25=2,p26=1,p27=0,p28=5,p29=5,p30=0,p31=0,p32=10,p33=2,p34=0,p35=0,p36=1,p37=1,p38=1,p39=1,p40=1,p41=1,p42=2,p43=5,p44=0,p45=5,p46=6,p47=0,p48=0,p49=10,p50=3,p51=0,p52=0,p53=1,p54=1,p55=1,p56=1,p57=1,p58=1,p59=9,p60=8,p61=0,p62=3,p63=9,p64=0,p65=0,p66=6,p67=8,p68=0,p69=0,p70=1,p71=1,p72=1,p73=1,p74=1,p75=1,p76=9,p77=1,p78=0,p79=3,p80=5,p81=0,p82=0,p83=6,p84=2,p85=0,p86=0,p87=1,p88=1,p89=1,p90=1,p91=1,p92=1,p93=9,p94=5,p95=0,p96=3,p97=6,p98=0,p99=0,p100=6,p101=3,p102=0,p103=0,p104=1,p105=1,p106=1,p107=1,p108=1,p109=1,p110=2,p111=8,p112=0,p113=2,p114=9,p115=0,p116=0,p117=6,p118=8,p119=0,p120=0,p121=1,p122=1,p123=1,p124=1,p125=1,p126=1,p127=2,p128=1,p129=0,p130=2,p131=5,p132=0,p133=0,p134=6,p135=2,p136=0,p137=0,p138=1,p139=1,p140=1,p141=1,p142=1,p143=1,p144=2,p145=5,p146=0,p147=2,p148=6,p149=0,p150=0,p151=6,p152=3,p153=0,p154=0,p155=0,p156=0,p157=1,p158=0,p159=1,p160=1,p161=1,p162=0,p163=1,p164=0,p165=1,p166=1,p167=0,p168=1,p169=1,p170=0,p171=1,p172=1,p173=1,p174=0,p175=1,p176=1,p177=1,p178=1,p179=0,p180=0,p181=1,p182=0,p183=1,p184=1,p185=1,p186=0,p187=1,p188=0,p189=1,p190=1,p191=0,p192=1,p193=1,p194=0,p195=1,p196=1,p197=1,p198=0,p199=1,p200=1,p201=1,p202=1,p203=0,p204=0,p205=0,p206=1,p207=1,p208=0,p209=1,p210=1,p211=1,p212=0,p213=1,p214=1,p215=1,p216=1,p217=0,p218=0,p219=1,p220=0,p221=1,p222=1,p223=1,p224=0,p225=1,p226=0,p227=1,p228=1,p229=0,p230=1,p231=1,p232=0,p233=1,p234=1,p235=1,p236=0,p237=1,p238=1,p239=1,p240=1,p241=0,p242=0,p243=0,p244=1,p245=1,p246=0,p247=1,p248=1,p249=1,p250=0,p251=1,p252=1,p253=1,p254=1,p255=0,p256=0,p257=1,p258=0,p259=1,p260=1,p261=1,p262=0,p263=1,p264=0,p265=1,p266=1,p267=0,p268=1,p269=1,p270=0,p271=1,p272=1,p273=1,p274=0,p275=1,p276=1,p277=1,p278=1,p279=0,p280=0,p281=1,p282=0,p283=1,p284=1,p285=1,p286=0,p287=1,p288=0,p289=1,p290=1,p291=0,p292=1,p293=1,p294=0,p295=1,p296=1,p297=1,p298=0,p299=1,p300=1,p301=1,p302=1,p303=0,p304=0,p305=0,p306=1,p307=1,p308=0,p309=1,p310=1,p311=1,p312=0,p313=1,p314=1,p315=1,p316=1,p317=0,p318=0,p319=1,p320=0,p321=1,p322=1,p323=1,p324=0,p325=1,p326=0,p327=1,p328=1,p329=0,p330=1,p331=1,p332=0,p333=1,p334=1,p335=1,p336=0,p337=1,p338=1,p339=1,p340=1,p341=0,p342=0,p343=0,p344=1,p345=1,p346=0,p347=1,p348=1,p349=1,p350=0,p351=1,p352=1,p353=1,p354=1,p355=0,p356=0,p357=1,p358=0,p359=1,p360=1,p361=1,p362=0,p363=1,p364=0,p365=1,p366=1,p367=0,p368=1,p369=1,p370=0,p371=1,p372=1,p373=1,p374=0,p375=1,p376=1,p377=1,p378=1,p379=0,p380=0,p381=1,p382=0,p383=1,p384=1,p385=1,p386=0,p387=1,p388=0,p389=1,p390=1,p391=0,p392=1,p393=1,p394=0,p395=1,p396=1,p397=1,p398=0,p399=1,p400=1,p401=1,p402=1,p403=0,p404=0,p405=0,p406=1,p407=1,p408=0,p409=1,p410=1,p411=1,p412=0,p413=1,p414=1,p415=1,p416=1,p417=0,p418=0,p419=1,p420=0,p421=1,p422=1,p423=1,p424=0,p425=1,p426=0,p427=1,p428=1,p429=0,p430=1,p431=1,p432=0,p433=1,p434=1,p435=1,p436=0,p437=1,p438=1,p439=1,p440=1,p441=0,p442=0,p443=0,p444=1,p445=1,p446=0,p447=1,p448=1,p449=1,p450=0,p451=1,p452=1,p453=1,p454=1,p455=0,p456=0,p457=1,p458=0,p459=1,p460=1,p461=1,p462=0,p463=1,p464=0,p465=1,p466=1,p467=0,p468=1,p469=1,p470=0,p471=1,p472=1,p473=1,p474=0,p475=1,p476=1,p477=1,p478=1,p479=0,p480=0,p481=1,p482=0,p483=1,p484=1,p485=1,p486=0,p487=1,p488=0,p489=1,p490=1,p491=0,p492=1,p493=1,p494=0,p495=1,p496=1,p497=1,p498=0,p499=1,p500=1,p501=1,p502=1,p503=0,p504=0,p505=0,p506=1,p507=1,p508=0,p509=1,p510=1,p511=1,p512=0,p513=1,p514=1,p515=1,p516=1,p517=0,p518=0,p519=1,p520=0,p521=1,p522=1,p523=1,p524=0,p525=1,p526=0,p527=1,p528=1,p529=0,p530=1,p531=1,p532=0,p533=1,p534=1,p535=1,p536=0,p537=1,p538=1,p539=1,p540=1,p541=0,p542=0,p543=0,p544=1,p545=1,p546=0,p547=1,p548=1,p549=1,p550=0,p551=1,p552=1,p553=1,p554=1,p555=0,p556=0,p557=1,p558=0,p559=1,p560=1,p561=1,p562=0,p563=1,p564=0,p565=1,p566=1,p567=0,p568=1,p569=1,p570=0,p571=1,p572=1,p573=1,p574=0,p575=1,p576=1,p577=1,p578=1,p579=0,p580=0,p581=1,p582=0,p583=1,p584=1,p585=1,p586=0,p587=1,p588=0,p589=1,p590=1,p591=0,p592=1,p593=1,p594=0,p595=1,p596=1,p597=1,p598=0,p599=1,p600=1,p601=1,p602=1,p603=0,p604=0,p605=0,p606=1,p607=1,p608=0,p609=1,p610=1,p611=1,p612=0,p613=1,p614=1,p615=1,p616=1,p617=0,p618=0,p619=1,p620=0,p621=1,p622=1,p623=1,p624=0,p625=1,p626=0,p627=1,p628=1,p629=0,p630=1,p631=1,p632=0,p633=1,p634=1,p635=1,p636=0,p637=1,p638=1,p639=1,p640=1,p641=0,p642=0,p643=0,p644=1,p645=1,p646=0,p647=1,p648=1,p649=1,p650=0,p651=1,p652=1,p653=1,p654=1,p655=0,p656=0,p657=1,p658=0,p659=1,p660=1,p661=1,p662=0,p663=1,p664=0,p665=1,p666=1,p667=0,p668=1,p669=1,p670=0,p671=1,p672=1,p673=1,p674=0,p675=1,p676=1,p677=1,p678=1,p679=0,p680=0,p681=1,p682=0,p683=1,p684=1,p685=1,p686=0,p687=1,p688=0,p689=1,p690=1,p691=0,p692=1,p693=1,p694=0,p695=1,p696=1,p697=1,p698=0,p699=1,p700=1,p701=1,p702=1,p703=0,p704=0,p705=0,p706=1,p707=1,p708=0,p709=1,p710=1,p711=1,p712=0,p713=1,p714=1,p715=1,p716=1,p717=0,p718=0,p719=1,p720=0,p721=1,p722=1,p723=1,p724=0,p725=1,p726=0,p727=1,p728=1,p729=0,p730=1,p731=1,p732=0,p733=1,p734=1,p735=1,p736=0,p737=1,p738=1,p739=1,p740=1,p741=0,p742=0,p743=0,p744=1,p745=1,p746=0,p747=1,p748=1,p749=1,p750=0,p751=1,p752=1,p753=1,p754=1,p755=0,p756=0,p757=1,p758=0,p759=1,p760=1,p761=1,p762=0,p763=1,p764=0,p765=1,p766=1,p767=0,p768=1,p769=1,p770=0,p771=1,p772=1,p773=1,p774=0,p775=1,p776=1,p777=1,p778=1,p779=0,p780=0,p781=1,p782=0,p783=1,p784=1,p785=1,p786=0,p787=1,p788=0,p789=1,p790=1,p791=0,p792=1,p793=1,p794=0,p795=1,p796=1,p797=1,p798=0,p799=1,p800=1,p801=1,p802=1,p803=0,p804=0,p805=0,p806=1,p807=1,p808=0,p809=1,p810=1,p811=1,p812=0,p813=1,p814=1,p815=1,p816=1,p817=0,p818=0,p819=1,p820=0,p821=1,p822=1,p823=1,p824=0,p825=1,p826=0,p827=1,p828=1,p829=0,p830=1,p831=1,p832=0,p833=1,p834=1,p835=1,p836=0,p837=1,p838=1,p839=1,p840=1,p841=0,p842=0,p843=0,p844=1,p845=1,p846=0,p847=1,p848=1,p849=1,p850=0,p851=1,p852=1,p853=1,p854=1,p855=0,p856=0,p857=1,p858=0,p859=1,p860=1,p861=1,p862=0,p863=1,p864=0,p865=1,p866=1,p867=0,p868=1,p869=1,p870=0,p871=1,p872=1,p873=1,p874=0,p875=1,p876=1,p877=1,p878=1,p879=0,p880=0,p881=1,p882=0,p883=1,p884=1,p885=1,p886=0,p887=1,p888=0,p889=1,p890=1,p891=0,p892=1,p893=1,p894=0,p895=1,p896=1,p897=1,p898=0,p899=1,p900=1,p901=1,p902=1,p903=0,p904=0,p905=0,p906=1,p907=1,p908=0,p909=1,p910=1,p911=1,p912=0,p913=1,p914=1,p915=1,p916=1,p917=0,p918=0,p919=1,p920=0,p921=1,p922=1,p923=1,p924=0,p925=1,p926=0,p927=1,p928=1,p929=0,p930=1,p931=1,p932=0,p933=1,p934=1,p935=1,p936=0,p937=1,p938=1,p939=1,p940=1,p941=0,p942=0,p943=0,p944=1,p945=1,p946=0,p947=1,p948=1,p949=1,p950=0,p951=1,p952=1,p953=1,p954=1,p955=0,p956=0,p957=1,p958=0,p959=1,p960=1,p961=1,p962=0,p963=1,p964=0,p965=1,p966=1,p967=0,p968=1,p969=1,p970=0,p971=1,p972=1,p973=1,p974=0,p975=1,p976=1,p977=1,p978=1,p979=0,p980=0,p981=1,p982=0,p983=1,p984=1,p985=1,p986=0,p987=1,p988=0,p989=1,p990=1,p991=0,p992=1,p993=1,p994=0,p995=1,p996=1,p997=1,p998=0,p999=1,p1000=1,p1001=1,p1002=1,p1003=0,p1004=0,p1005=0,p1006=1,p1007=1,p1008=0,p1009=1,p1010=1,p1011=1,p1012=0,p1013=1,p1014=1,p1015=1,p1016=1,p1017=0,p1018=0,p1019=1,p1020=0,p1021=1,p1022=1,p1023=1,p1024=0,p1025=1,p1026=0,p1027=1,p1028=1,p1029=0,p1030=1,p1031=1,p1032=0,p1033=1,p1034=1,p1035=1,p1036=0,p1037=1,p1038=1,p1039=1,p1040=1,p1041=0,p1042=0,p1043=0,p1044=1,p1045=1,p1046=0,p1047=1,p1048=1,p1049=1,p1050=0,p1051=1,p1052=1,p1053=1,p1054=1;
reg [11:0] f0,f1,f2,f3,f4,f5,f6,f7,f8,f9,f10,f11,f12,f13,f14,f15,f16,f17,f18,f19,f20,f21,f22,f23,f24,f25,f26,f27,f28,f29,f30,f31,f32,f33,f34,f35,f36,f37,f38,f39,f40,f41,f42,f43,f44,f45,f46,f47,f48,f49,f50,f51,f52,f53,f54,f55,f56,f57,f58,f59,f60,f61,f62,f63,f64,f65,f66,f67,f68,f69,f70,f71,f72,f73,f74,f75,f76,f77,f78,f79,f80,f81,f82,f83,f84,f85,f86,f87,f88,f89,f90,f91,f92,f93,f94,f95,f96,f97,f98,f99,f100,f101,f102,f103,f104,f105,f106,f107,f108,f109,f110,f111,f112,f113,f114,f115,f116,f117,f118,f119,f120,f121,f122,f123,f124,f125,f126,f127,f128,f129,f130,f131,f132,f133,f134,f135,f136,f137,f138,f139,f140,f141,f142,f143,f144,f145,f146,f147,f148,f149,f150,f151,f152,f153,f154,f155,f156,f157,f158,f159,f160,f161,f162,f163,f164,f165,f166,f167,f168,f169,f170,f171,f172,f173,f174,f175,f176,f177,f178,f179,f180,f181,f182,f183,f184,f185,f186,f187,f188,f189,f190,f191,f192,f193,f194,f195,f196,f197,f198,f199,f200,f201,f202,f203,f204,f205,f206,f207,f208,f209,f210,f211,f212,f213,f214,f215,f216,f217,f218,f219,f220,f221,f222,f223,f224,f225,f226,f227,f228,f229,f230,f231,f232,f233,f234,f235,f236,f237,f238,f239,f240,f241,f242,f243,f244,f245,f246,f247,f248,f249,f250,f251,f252,f253,f254,f255,f256,f257,f258,f259,f260,f261,f262,f263,f264,f265,f266,f267,f268,f269,f270,f271,f272,f273,f274,f275,f276,f277,f278,f279,f280,f281,f282,f283,f284,f285,f286,f287,f288,f289,f290,f291,f292,f293,f294,f295,f296,f297,f298,f299,f300,f301,f302,f303,f304,f305,f306,f307,f308,f309,f310,f311,f312,f313,f314,f315,f316,f317,f318,f319,f320,f321,f322,f323,f324,f325,f326,f327,f328,f329,f330,f331,f332,f333,f334,f335,f336,f337,f338,f339,f340,f341,f342,f343,f344,f345,f346,f347,f348,f349,f350,f351,f352,f353,f354,f355,f356,f357,f358,f359,f360,f361,f362,f363,f364,f365,f366,f367,f368,f369,f370,f371,f372,f373,f374,f375,f376,f377,f378,f379,f380,f381,f382,f383,f384,f385,f386,f387,f388,f389,f390,f391,f392,f393,f394,f395,f396,f397,f398,f399,f400,f401,f402,f403,f404,f405,f406,f407,f408,f409,f410,f411,f412,f413,f414,f415,f416,f417,f418,f419,f420,f421,f422,f423,f424,f425,f426,f427,f428,f429,f430,f431,f432,f433,f434,f435,f436,f437,f438,f439,f440,f441,f442,f443,f444,f445,f446,f447,f448,f449,f450,f451,f452,f453,f454,f455,f456,f457,f458,f459,f460,f461,f462,f463,f464,f465,f466,f467,f468,f469,f470,f471,f472,f473,f474,f475,f476,f477,f478,f479,f480,f481,f482,f483,f484,f485,f486,f487,f488,f489,f490,f491,f492,f493,f494,f495,f496,f497,f498,f499,f500,f501,f502,f503,f504,f505,f506,f507,f508,f509,f510,f511,f512,f513,f514,f515,f516,f517,f518,f519,f520,f521,f522,f523,f524,f525,f526,f527,f528,f529,f530,f531,f532,f533,f534,f535,f536,f537,f538,f539,f540,f541,f542,f543,f544,f545,f546,f547,f548,f549,f550,f551,f552,f553,f554,f555,f556,f557,f558,f559,f560,f561,f562,f563,f564,f565,f566,f567,f568,f569,f570,f571,f572,f573,f574,f575,f576,f577,f578,f579,f580,f581,f582,f583,f584,f585,f586,f587,f588,f589,f590,f591,f592,f593,f594,f595,f596,f597,f598,f599,f600,f601,f602,f603,f604,f605,f606,f607,f608,f609,f610,f611,f612,f613,f614,f615,f616,f617,f618,f619,f620,f621,f622,f623,f624,f625,f626,f627,f628,f629,f630,f631,f632,f633,f634,f635,f636,f637,f638,f639,f640,f641,f642,f643,f644,f645,f646,f647,f648,f649,f650,f651,f652,f653,f654,f655,f656,f657,f658,f659,f660,f661,f662,f663,f664,f665,f666,f667,f668,f669,f670,f671,f672,f673,f674,f675,f676,f677,f678,f679,f680,f681,f682,f683,f684,f685,f686,f687,f688,f689,f690,f691,f692,f693,f694,f695,f696,f697,f698,f699,f700,f701,f702,f703,f704,f705,f706,f707,f708,f709,f710,f711,f712,f713,f714,f715,f716,f717,f718,f719,f720,f721,f722,f723,f724,f725,f726,f727,f728,f729,f730,f731,f732,f733,f734,f735,f736,f737,f738,f739,f740,f741,f742,f743,f744,f745,f746,f747,f748,f749,f750,f751,f752,f753,f754,f755,f756,f757,f758,f759,f760,f761,f762,f763,f764,f765,f766,f767,f768,f769,f770,f771,f772,f773,f774,f775,f776,f777,f778,f779,f780,f781,f782,f783,f784,f785,f786,f787,f788,f789,f790,f791,f792,f793,f794,f795,f796,f797,f798,f799,f800,f801,f802,f803,f804,f805,f806,f807,f808,f809,f810,f811,f812,f813,f814,f815,f816,f817,f818,f819,f820,f821,f822,f823,f824,f825,f826,f827,f828,f829,f830,f831,f832,f833,f834,f835,f836,f837,f838,f839,f840,f841,f842,f843,f844,f845,f846,f847,f848,f849,f850,f851,f852,f853,f854,f855,f856,f857,f858,f859,f860,f861,f862,f863,f864,f865,f866,f867,f868,f869,f870,f871,f872,f873,f874,f875,f876,f877,f878,f879,f880,f881,f882,f883,f884,f885,f886,f887,f888,f889,f890,f891,f892,f893,f894,f895,f896,f897,f898,f899,f900,f901,f902,f903,f904,f905,f906,f907,f908,f909,f910,f911,f912,f913,f914,f915,f916,f917,f918,f919,f920,f921,f922,f923,f924,f925,f926,f927,f928,f929,f930,f931,f932,f933,f934,f935,f936,f937,f938,f939,f940,f941,f942,f943,f944,f945,f946,f947,f948,f949,f950,f951,f952,f953,f954,f955,f956,f957,f958,f959,f960,f961,f962,f963,f964,f965,f966,f967,f968,f969,f970,f971,f972,f973,f974,f975,f976,f977,f978,f979,f980,f981,f982,f983,f984,f985,f986,f987,f988,f989,f990,f991,f992,f993,f994,f995,f996,f997,f998,f999,f1000,f1001,f1002,f1003,f1004,f1005,f1006,f1007,f1008,f1009,f1010,f1011,f1012,f1013,f1014,f1015,f1016,f1017,f1018,f1019,f1020,f1021,f1022,f1023,f1024,f1025,f1026,f1027,f1028,f1029,f1030,f1031,f1032,f1033,f1034,f1035,f1036,f1037,f1038,f1039,f1040,f1041,f1042,f1043,f1044,f1045,f1046,f1047,f1048,f1049,f1050,f1051,f1052,f1053,f1054,f1055,f1056,f1057,f1058,f1059,f1060,f1061,f1062,f1063,f1064,f1065,f1066,f1067,f1068,f1069,f1070,f1071,f1072,f1073,f1074,f1075,f1076,f1077,f1078,f1079,f1080,f1081,f1082,f1083,f1084,f1085,f1086,f1087,f1088,f1089,f1090,f1091,f1092,f1093,f1094,f1095,f1096,f1097,f1098,f1099,f1100,f1101,f1102,f1103,f1104,f1105,f1106,f1107,f1108,f1109,f1110,f1111,f1112,f1113,f1114,f1115,f1116,f1117;
reg [11:0] tf;
reg [11:0] tc;
reg [1:0] clk_div; // 2位寄存器用于实现时钟分频
reg [47:0] counter1=1;
always @(posedge clk) begin
    if(clk_div < 2'b11)
        clk_div <= clk_div + 1; // 计数器自增
    else
        clk_div <= 2'b00; // 重置计数器
end

// 使用clk_div来控制某些逻辑的触发条件
always @(posedge clk) begin
    if (clk_div == 2'b11) begin
        f0 = 4095;
        f0 = (f0 >= `INH(p0)) ? `INH(p0) : f0;
        f0 = (f0 > p2) ? p2 : f0;
        f0 = (f0 > p19) ? p19 : f0;
        f0 = (f0 > p36) ? p36 : f0;
        f0 = (f0 > p53) ? p53 : f0;
        f0 = (f0 > p70) ? p70 : f0;
        f0 = (f0 > p87) ? p87 : f0;
        f0 = (f0 > p104) ? p104 : f0;
        f0 = (f0 > p121) ? p121 : f0;
        f0 = (f0 > p138) ? p138 : f0;
        f1 = 4095;
        f1 = (f1 > p1) ? p1 : f1;
        f1 = (f1 >= `INH(p7)) ? `INH(p7) : f1;
        f1 = (f1 >= `INH(p24)) ? `INH(p24) : f1;
        f1 = (f1 >= `INH(p41)) ? `INH(p41) : f1;
        f1 = (f1 >= `INH(p58)) ? `INH(p58) : f1;
        f1 = (f1 >= `INH(p75)) ? `INH(p75) : f1;
        f1 = (f1 >= `INH(p92)) ? `INH(p92) : f1;
        f1 = (f1 >= `INH(p109)) ? `INH(p109) : f1;
        f1 = (f1 >= `INH(p126)) ? `INH(p126) : f1;
        f1 = (f1 >= `INH(p143)) ? `INH(p143) : f1;
        f2 = 4095;
        f2 = (f2 >= `INH(p157)) ? `INH(p157) : f2;
        f2 = (f2 > p160) ? p160 : f2;
        f3 = 4095;
        f3 = (f3 >= `INH(p181)) ? `INH(p181) : f3;
        f3 = (f3 > p184) ? p184 : f3;
        f4 = 4095;
        f4 = (f4 > p203) ? p203 : f4;
        f4 = (f4 >= `INH(p206)) ? `INH(p206) : f4;
        f5 = 4095;
        f5 = (f5 >= `INH(p219)) ? `INH(p219) : f5;
        f5 = (f5 > p222) ? p222 : f5;
        f6 = 4095;
        f6 = (f6 > p241) ? p241 : f6;
        f6 = (f6 >= `INH(p244)) ? `INH(p244) : f6;
        f7 = 4095;
        f7 = (f7 >= `INH(p257)) ? `INH(p257) : f7;
        f7 = (f7 > p260) ? p260 : f7;
        f8 = 4095;
        f8 = (f8 >= `INH(p281)) ? `INH(p281) : f8;
        f8 = (f8 > p284) ? p284 : f8;
        f9 = 4095;
        f9 = (f9 > p303) ? p303 : f9;
        f9 = (f9 >= `INH(p306)) ? `INH(p306) : f9;
        f10 = 4095;
        f10 = (f10 >= `INH(p319)) ? `INH(p319) : f10;
        f10 = (f10 > p322) ? p322 : f10;
        f11 = 4095;
        f11 = (f11 > p341) ? p341 : f11;
        f11 = (f11 >= `INH(p344)) ? `INH(p344) : f11;
        f12 = 4095;
        f12 = (f12 >= `INH(p357)) ? `INH(p357) : f12;
        f12 = (f12 > p360) ? p360 : f12;
        f13 = 4095;
        f13 = (f13 >= `INH(p381)) ? `INH(p381) : f13;
        f13 = (f13 > p384) ? p384 : f13;
        f14 = 4095;
        f14 = (f14 > p403) ? p403 : f14;
        f14 = (f14 >= `INH(p406)) ? `INH(p406) : f14;
        f15 = 4095;
        f15 = (f15 >= `INH(p419)) ? `INH(p419) : f15;
        f15 = (f15 > p422) ? p422 : f15;
        f16 = 4095;
        f16 = (f16 > p441) ? p441 : f16;
        f16 = (f16 >= `INH(p444)) ? `INH(p444) : f16;
        f17 = 4095;
        f17 = (f17 >= `INH(p457)) ? `INH(p457) : f17;
        f17 = (f17 > p460) ? p460 : f17;
        f18 = 4095;
        f18 = (f18 >= `INH(p481)) ? `INH(p481) : f18;
        f18 = (f18 > p484) ? p484 : f18;
        f19 = 4095;
        f19 = (f19 > p503) ? p503 : f19;
        f19 = (f19 >= `INH(p506)) ? `INH(p506) : f19;
        f20 = 4095;
        f20 = (f20 >= `INH(p519)) ? `INH(p519) : f20;
        f20 = (f20 > p522) ? p522 : f20;
        f21 = 4095;
        f21 = (f21 > p541) ? p541 : f21;
        f21 = (f21 >= `INH(p544)) ? `INH(p544) : f21;
        f22 = 4095;
        f22 = (f22 >= `INH(p557)) ? `INH(p557) : f22;
        f22 = (f22 > p560) ? p560 : f22;
        f23 = 4095;
        f23 = (f23 >= `INH(p581)) ? `INH(p581) : f23;
        f23 = (f23 > p584) ? p584 : f23;
        f24 = 4095;
        f24 = (f24 > p603) ? p603 : f24;
        f24 = (f24 >= `INH(p606)) ? `INH(p606) : f24;
        f25 = 4095;
        f25 = (f25 >= `INH(p619)) ? `INH(p619) : f25;
        f25 = (f25 > p622) ? p622 : f25;
        f26 = 4095;
        f26 = (f26 > p641) ? p641 : f26;
        f26 = (f26 >= `INH(p644)) ? `INH(p644) : f26;
        f27 = 4095;
        f27 = (f27 >= `INH(p657)) ? `INH(p657) : f27;
        f27 = (f27 > p660) ? p660 : f27;
        f28 = 4095;
        f28 = (f28 >= `INH(p681)) ? `INH(p681) : f28;
        f28 = (f28 > p684) ? p684 : f28;
        f29 = 4095;
        f29 = (f29 > p703) ? p703 : f29;
        f29 = (f29 >= `INH(p706)) ? `INH(p706) : f29;
        f30 = 4095;
        f30 = (f30 >= `INH(p719)) ? `INH(p719) : f30;
        f30 = (f30 > p722) ? p722 : f30;
        f31 = 4095;
        f31 = (f31 > p741) ? p741 : f31;
        f31 = (f31 >= `INH(p744)) ? `INH(p744) : f31;
        f32 = 4095;
        f32 = (f32 >= `INH(p757)) ? `INH(p757) : f32;
        f32 = (f32 > p760) ? p760 : f32;
        f33 = 4095;
        f33 = (f33 >= `INH(p781)) ? `INH(p781) : f33;
        f33 = (f33 > p784) ? p784 : f33;
        f34 = 4095;
        f34 = (f34 > p803) ? p803 : f34;
        f34 = (f34 >= `INH(p806)) ? `INH(p806) : f34;
        f35 = 4095;
        f35 = (f35 >= `INH(p819)) ? `INH(p819) : f35;
        f35 = (f35 > p822) ? p822 : f35;
        f36 = 4095;
        f36 = (f36 > p841) ? p841 : f36;
        f36 = (f36 >= `INH(p844)) ? `INH(p844) : f36;
        f37 = 4095;
        f37 = (f37 >= `INH(p857)) ? `INH(p857) : f37;
        f37 = (f37 > p860) ? p860 : f37;
        f38 = 4095;
        f38 = (f38 >= `INH(p881)) ? `INH(p881) : f38;
        f38 = (f38 > p884) ? p884 : f38;
        f39 = 4095;
        f39 = (f39 > p903) ? p903 : f39;
        f39 = (f39 >= `INH(p906)) ? `INH(p906) : f39;
        f40 = 4095;
        f40 = (f40 >= `INH(p919)) ? `INH(p919) : f40;
        f40 = (f40 > p922) ? p922 : f40;
        f41 = 4095;
        f41 = (f41 > p941) ? p941 : f41;
        f41 = (f41 >= `INH(p944)) ? `INH(p944) : f41;
        f42 = 4095;
        f42 = (f42 >= `INH(p957)) ? `INH(p957) : f42;
        f42 = (f42 > p960) ? p960 : f42;
        f43 = 4095;
        f43 = (f43 >= `INH(p981)) ? `INH(p981) : f43;
        f43 = (f43 > p984) ? p984 : f43;
        f44 = 4095;
        f44 = (f44 > p1003) ? p1003 : f44;
        f44 = (f44 >= `INH(p1006)) ? `INH(p1006) : f44;
        f45 = 4095;
        f45 = (f45 >= `INH(p1019)) ? `INH(p1019) : f45;
        f45 = (f45 > p1022) ? p1022 : f45;
        f46 = 4095;
        f46 = (f46 > p1041) ? p1041 : f46;
        f46 = (f46 >= `INH(p1044)) ? `INH(p1044) : f46;
        f47 = 4095;
        f47 = (f47 >= `INH(p156)) ? `INH(p156) : f47;
        f47 = (f47 >= `INH(p157)) ? `INH(p157) : f47;
        f47 = (f47 > p161) ? p161 : f47;
        f48 = 4095;
        f48 = (f48 > p155) ? p155 : f48;
        f48 = (f48 >= `INH(p161)) ? `INH(p161) : f48;
        f49 = 4095;
        f49 = (f49 > p159) ? p159 : f49;
        f49 = (f49 >= `INH(p161)) ? `INH(p161) : f49;
        f50 = 4095;
        f50 = (f50 >= p156/2) ? p156/2 : f50;
        f50 = (f50 >= `INH(p160)) ? `INH(p160) : f50;
        f51 = 4095;
        f51 = (f51 >= `INH(p160)) ? `INH(p160) : f51;
        f51 = (f51 > p163) ? p163 : f51;
        f52 = 4095;
        f52 = (f52 > p156) ? p156 : f52;
        f52 = (f52 >= `INH(p163)) ? `INH(p163) : f52;
        f52 = (f52 > p165) ? p165 : f52;
        f53 = 4095;
        f53 = (f53 >= `INH(p163)) ? `INH(p163) : f53;
        f53 = (f53 > p166) ? p166 : f53;
        f54 = 4095;
        f54 = (f54 > p155) ? p155 : f54;
        f54 = (f54 >= `INH(p165)) ? `INH(p165) : f54;
        f54 = (f54 >= `INH(p166)) ? `INH(p166) : f54;
        f55 = 4095;
        f55 = (f55 > p155) ? p155 : f55;
        f55 = (f55 >= `INH(p164)) ? `INH(p164) : f55;
        f55 = (f55 >= `INH(p166)) ? `INH(p166) : f55;
        f56 = 4095;
        f56 = (f56 >= `INH(p166)) ? `INH(p166) : f56;
        f56 = (f56 > p168) ? p168 : f56;
        f57 = 4095;
        f57 = (f57 > p162) ? p162 : f57;
        f57 = (f57 >= `INH(p168)) ? `INH(p168) : f57;
        f58 = 4095;
        f58 = (f58 >= `INH(p168)) ? `INH(p168) : f58;
        f58 = (f58 > p169) ? p169 : f58;
        f59 = 4095;
        f59 = (f59 > p167) ? p167 : f59;
        f59 = (f59 >= `INH(p169)) ? `INH(p169) : f59;
        f60 = 4095;
        f60 = (f60 > p157) ? p157 : f60;
        f60 = (f60 > p164) ? p164 : f60;
        f60 = (f60 >= `INH(p165)) ? `INH(p165) : f60;
        f60 = (f60 >= `INH(p169)) ? `INH(p169) : f60;
        f61 = 4095;
        f61 = (f61 > p157) ? p157 : f61;
        f61 = (f61 >= `INH(p164)) ? `INH(p164) : f61;
        f61 = (f61 >= `INH(p169)) ? `INH(p169) : f61;
        f62 = 4095;
        f62 = (f62 > p8) ? p8 : f62;
        f62 = (f62 >= `INH(p171)) ? `INH(p171) : f62;
        f63 = 4095;
        f63 = (f63 > p170) ? p170 : f63;
        f63 = (f63 >= `INH(p172)) ? `INH(p172) : f63;
        f64 = 4095;
        f64 = (f64 >= `INH(p8)) ? `INH(p8) : f64;
        f64 = (f64 >= `INH(p171)) ? `INH(p171) : f64;
        f64 = (f64 > p172) ? p172 : f64;
        f65 = 4095;
        f65 = (f65 >= `INH(p170)) ? `INH(p170) : f65;
        f65 = (f65 >= `INH(p172)) ? `INH(p172) : f65;
        f65 = (f65 > p173) ? p173 : f65;
        f66 = 4095;
        f66 = (f66 > p9) ? p9 : f66;
        f66 = (f66 >= `INH(p175)) ? `INH(p175) : f66;
        f67 = 4095;
        f67 = (f67 > p174) ? p174 : f67;
        f67 = (f67 >= `INH(p176)) ? `INH(p176) : f67;
        f68 = 4095;
        f68 = (f68 >= `INH(p9)) ? `INH(p9) : f68;
        f68 = (f68 >= `INH(p175)) ? `INH(p175) : f68;
        f68 = (f68 > p176) ? p176 : f68;
        f69 = 4095;
        f69 = (f69 >= `INH(p174)) ? `INH(p174) : f69;
        f69 = (f69 >= `INH(p176)) ? `INH(p176) : f69;
        f69 = (f69 > p177) ? p177 : f69;
        f70 = 4095;
        f70 = (f70 >= `INH(p2)) ? `INH(p2) : f70;
        f70 = (f70 > p171) ? p171 : f70;
        f70 = (f70 > p175) ? p175 : f70;
        f71 = 4095;
        f71 = (f71 > p157) ? p157 : f71;
        f71 = (f71 >= `INH(p173)) ? `INH(p173) : f71;
        f71 = (f71 >= `INH(p177)) ? `INH(p177) : f71;
        f72 = 4095;
        f72 = (f72 > p158) ? p158 : f72;
        f72 = (f72 >= `INH(p178)) ? `INH(p178) : f72;
        f73 = 4095;
        f73 = (f73 > p10) ? p10 : f73;
        f73 = (f73 >= `INH(p159)) ? `INH(p159) : f73;
        f74 = 4095;
        f74 = (f74 >= `INH(p10)) ? `INH(p10) : f74;
        f74 = (f74 >= `INH(p159)) ? `INH(p159) : f74;
        f74 = (f74 > p178) ? p178 : f74;
        f75 = 4095;
        f75 = (f75 > p3) ? p3 : f75;
        f75 = (f75 >= `INH(p158)) ? `INH(p158) : f75;
        f75 = (f75 >= `INH(p178)) ? `INH(p178) : f75;
        f76 = 4095;
        f76 = (f76 >= `INH(p180)) ? `INH(p180) : f76;
        f76 = (f76 >= `INH(p181)) ? `INH(p181) : f76;
        f76 = (f76 > p185) ? p185 : f76;
        f77 = 4095;
        f77 = (f77 > p179) ? p179 : f77;
        f77 = (f77 >= `INH(p185)) ? `INH(p185) : f77;
        f78 = 4095;
        f78 = (f78 > p183) ? p183 : f78;
        f78 = (f78 >= `INH(p185)) ? `INH(p185) : f78;
        f79 = 4095;
        f79 = (f79 >= p180/2) ? p180/2 : f79;
        f79 = (f79 >= `INH(p184)) ? `INH(p184) : f79;
        f80 = 4095;
        f80 = (f80 >= `INH(p184)) ? `INH(p184) : f80;
        f80 = (f80 > p187) ? p187 : f80;
        f81 = 4095;
        f81 = (f81 > p180) ? p180 : f81;
        f81 = (f81 >= `INH(p187)) ? `INH(p187) : f81;
        f81 = (f81 > p189) ? p189 : f81;
        f82 = 4095;
        f82 = (f82 >= `INH(p187)) ? `INH(p187) : f82;
        f82 = (f82 > p190) ? p190 : f82;
        f83 = 4095;
        f83 = (f83 > p179) ? p179 : f83;
        f83 = (f83 >= `INH(p189)) ? `INH(p189) : f83;
        f83 = (f83 >= `INH(p190)) ? `INH(p190) : f83;
        f84 = 4095;
        f84 = (f84 > p179) ? p179 : f84;
        f84 = (f84 >= `INH(p188)) ? `INH(p188) : f84;
        f84 = (f84 >= `INH(p190)) ? `INH(p190) : f84;
        f85 = 4095;
        f85 = (f85 >= `INH(p190)) ? `INH(p190) : f85;
        f85 = (f85 > p192) ? p192 : f85;
        f86 = 4095;
        f86 = (f86 > p186) ? p186 : f86;
        f86 = (f86 >= `INH(p192)) ? `INH(p192) : f86;
        f87 = 4095;
        f87 = (f87 >= `INH(p192)) ? `INH(p192) : f87;
        f87 = (f87 > p193) ? p193 : f87;
        f88 = 4095;
        f88 = (f88 > p191) ? p191 : f88;
        f88 = (f88 >= `INH(p193)) ? `INH(p193) : f88;
        f89 = 4095;
        f89 = (f89 > p181) ? p181 : f89;
        f89 = (f89 > p188) ? p188 : f89;
        f89 = (f89 >= `INH(p189)) ? `INH(p189) : f89;
        f89 = (f89 >= `INH(p193)) ? `INH(p193) : f89;
        f90 = 4095;
        f90 = (f90 > p181) ? p181 : f90;
        f90 = (f90 >= `INH(p188)) ? `INH(p188) : f90;
        f90 = (f90 >= `INH(p193)) ? `INH(p193) : f90;
        f91 = 4095;
        f91 = (f91 > p11) ? p11 : f91;
        f91 = (f91 >= `INH(p195)) ? `INH(p195) : f91;
        f92 = 4095;
        f92 = (f92 > p194) ? p194 : f92;
        f92 = (f92 >= `INH(p196)) ? `INH(p196) : f92;
        f93 = 4095;
        f93 = (f93 >= `INH(p11)) ? `INH(p11) : f93;
        f93 = (f93 >= `INH(p195)) ? `INH(p195) : f93;
        f93 = (f93 > p196) ? p196 : f93;
        f94 = 4095;
        f94 = (f94 >= `INH(p194)) ? `INH(p194) : f94;
        f94 = (f94 >= `INH(p196)) ? `INH(p196) : f94;
        f94 = (f94 > p197) ? p197 : f94;
        f95 = 4095;
        f95 = (f95 > p12) ? p12 : f95;
        f95 = (f95 >= `INH(p199)) ? `INH(p199) : f95;
        f96 = 4095;
        f96 = (f96 > p198) ? p198 : f96;
        f96 = (f96 >= `INH(p200)) ? `INH(p200) : f96;
        f97 = 4095;
        f97 = (f97 >= `INH(p12)) ? `INH(p12) : f97;
        f97 = (f97 >= `INH(p199)) ? `INH(p199) : f97;
        f97 = (f97 > p200) ? p200 : f97;
        f98 = 4095;
        f98 = (f98 >= `INH(p198)) ? `INH(p198) : f98;
        f98 = (f98 >= `INH(p200)) ? `INH(p200) : f98;
        f98 = (f98 > p201) ? p201 : f98;
        f99 = 4095;
        f99 = (f99 >= `INH(p3)) ? `INH(p3) : f99;
        f99 = (f99 > p195) ? p195 : f99;
        f99 = (f99 > p199) ? p199 : f99;
        f100 = 4095;
        f100 = (f100 > p181) ? p181 : f100;
        f100 = (f100 >= `INH(p197)) ? `INH(p197) : f100;
        f100 = (f100 >= `INH(p201)) ? `INH(p201) : f100;
        f101 = 4095;
        f101 = (f101 > p182) ? p182 : f101;
        f101 = (f101 >= `INH(p202)) ? `INH(p202) : f101;
        f102 = 4095;
        f102 = (f102 > p13) ? p13 : f102;
        f102 = (f102 >= `INH(p183)) ? `INH(p183) : f102;
        f103 = 4095;
        f103 = (f103 >= `INH(p13)) ? `INH(p13) : f103;
        f103 = (f103 >= `INH(p183)) ? `INH(p183) : f103;
        f103 = (f103 > p202) ? p202 : f103;
        f104 = 4095;
        f104 = (f104 > p4) ? p4 : f104;
        f104 = (f104 >= `INH(p182)) ? `INH(p182) : f104;
        f104 = (f104 >= `INH(p202)) ? `INH(p202) : f104;
        f105 = 4095;
        f105 = (f105 > p204) ? p204 : f105;
        f105 = (f105 >= `INH(p206)) ? `INH(p206) : f105;
        f106 = 4095;
        f106 = (f106 >= `INH(p203)) ? `INH(p203) : f106;
        f106 = (f106 >= `INH(p204)) ? `INH(p204) : f106;
        f106 = (f106 >= `INH(p206)) ? `INH(p206) : f106;
        f106 = (f106 > p207) ? p207 : f106;
        f107 = 4095;
        f107 = (f107 > p10) ? p10 : f107;
        f107 = (f107 >= `INH(p209)) ? `INH(p209) : f107;
        f108 = 4095;
        f108 = (f108 > p208) ? p208 : f108;
        f108 = (f108 >= `INH(p210)) ? `INH(p210) : f108;
        f109 = 4095;
        f109 = (f109 >= `INH(p10)) ? `INH(p10) : f109;
        f109 = (f109 >= `INH(p209)) ? `INH(p209) : f109;
        f109 = (f109 > p210) ? p210 : f109;
        f110 = 4095;
        f110 = (f110 >= `INH(p208)) ? `INH(p208) : f110;
        f110 = (f110 >= `INH(p210)) ? `INH(p210) : f110;
        f110 = (f110 > p211) ? p211 : f110;
        f111 = 4095;
        f111 = (f111 > p13) ? p13 : f111;
        f111 = (f111 >= `INH(p213)) ? `INH(p213) : f111;
        f112 = 4095;
        f112 = (f112 > p212) ? p212 : f112;
        f112 = (f112 >= `INH(p214)) ? `INH(p214) : f112;
        f113 = 4095;
        f113 = (f113 >= `INH(p13)) ? `INH(p13) : f113;
        f113 = (f113 >= `INH(p213)) ? `INH(p213) : f113;
        f113 = (f113 > p214) ? p214 : f113;
        f114 = 4095;
        f114 = (f114 >= `INH(p212)) ? `INH(p212) : f114;
        f114 = (f114 >= `INH(p214)) ? `INH(p214) : f114;
        f114 = (f114 > p215) ? p215 : f114;
        f115 = 4095;
        f115 = (f115 >= `INH(p4)) ? `INH(p4) : f115;
        f115 = (f115 > p209) ? p209 : f115;
        f115 = (f115 > p213) ? p213 : f115;
        f116 = 4095;
        f116 = (f116 > p206) ? p206 : f116;
        f116 = (f116 >= `INH(p211)) ? `INH(p211) : f116;
        f116 = (f116 >= `INH(p215)) ? `INH(p215) : f116;
        f117 = 4095;
        f117 = (f117 > p205) ? p205 : f117;
        f117 = (f117 >= `INH(p216)) ? `INH(p216) : f117;
        f118 = 4095;
        f118 = (f118 > p14) ? p14 : f118;
        f118 = (f118 >= `INH(p207)) ? `INH(p207) : f118;
        f119 = 4095;
        f119 = (f119 >= `INH(p14)) ? `INH(p14) : f119;
        f119 = (f119 >= `INH(p207)) ? `INH(p207) : f119;
        f119 = (f119 > p216) ? p216 : f119;
        f120 = 4095;
        f120 = (f120 > p5) ? p5 : f120;
        f120 = (f120 >= `INH(p205)) ? `INH(p205) : f120;
        f120 = (f120 >= `INH(p216)) ? `INH(p216) : f120;
        f121 = 4095;
        f121 = (f121 >= `INH(p218)) ? `INH(p218) : f121;
        f121 = (f121 >= `INH(p219)) ? `INH(p219) : f121;
        f121 = (f121 > p223) ? p223 : f121;
        f122 = 4095;
        f122 = (f122 > p217) ? p217 : f122;
        f122 = (f122 >= `INH(p223)) ? `INH(p223) : f122;
        f123 = 4095;
        f123 = (f123 > p221) ? p221 : f123;
        f123 = (f123 >= `INH(p223)) ? `INH(p223) : f123;
        f124 = 4095;
        f124 = (f124 >= p218/2) ? p218/2 : f124;
        f124 = (f124 >= `INH(p222)) ? `INH(p222) : f124;
        f125 = 4095;
        f125 = (f125 >= `INH(p222)) ? `INH(p222) : f125;
        f125 = (f125 > p225) ? p225 : f125;
        f126 = 4095;
        f126 = (f126 > p218) ? p218 : f126;
        f126 = (f126 >= `INH(p225)) ? `INH(p225) : f126;
        f126 = (f126 > p227) ? p227 : f126;
        f127 = 4095;
        f127 = (f127 >= `INH(p225)) ? `INH(p225) : f127;
        f127 = (f127 > p228) ? p228 : f127;
        f128 = 4095;
        f128 = (f128 > p217) ? p217 : f128;
        f128 = (f128 >= `INH(p227)) ? `INH(p227) : f128;
        f128 = (f128 >= `INH(p228)) ? `INH(p228) : f128;
        f129 = 4095;
        f129 = (f129 > p217) ? p217 : f129;
        f129 = (f129 >= `INH(p226)) ? `INH(p226) : f129;
        f129 = (f129 >= `INH(p228)) ? `INH(p228) : f129;
        f130 = 4095;
        f130 = (f130 >= `INH(p228)) ? `INH(p228) : f130;
        f130 = (f130 > p230) ? p230 : f130;
        f131 = 4095;
        f131 = (f131 > p224) ? p224 : f131;
        f131 = (f131 >= `INH(p230)) ? `INH(p230) : f131;
        f132 = 4095;
        f132 = (f132 >= `INH(p230)) ? `INH(p230) : f132;
        f132 = (f132 > p231) ? p231 : f132;
        f133 = 4095;
        f133 = (f133 > p229) ? p229 : f133;
        f133 = (f133 >= `INH(p231)) ? `INH(p231) : f133;
        f134 = 4095;
        f134 = (f134 > p219) ? p219 : f134;
        f134 = (f134 > p226) ? p226 : f134;
        f134 = (f134 >= `INH(p227)) ? `INH(p227) : f134;
        f134 = (f134 >= `INH(p231)) ? `INH(p231) : f134;
        f135 = 4095;
        f135 = (f135 > p219) ? p219 : f135;
        f135 = (f135 >= `INH(p226)) ? `INH(p226) : f135;
        f135 = (f135 >= `INH(p231)) ? `INH(p231) : f135;
        f136 = 4095;
        f136 = (f136 > p15) ? p15 : f136;
        f136 = (f136 >= `INH(p233)) ? `INH(p233) : f136;
        f137 = 4095;
        f137 = (f137 > p232) ? p232 : f137;
        f137 = (f137 >= `INH(p234)) ? `INH(p234) : f137;
        f138 = 4095;
        f138 = (f138 >= `INH(p15)) ? `INH(p15) : f138;
        f138 = (f138 >= `INH(p233)) ? `INH(p233) : f138;
        f138 = (f138 > p234) ? p234 : f138;
        f139 = 4095;
        f139 = (f139 >= `INH(p232)) ? `INH(p232) : f139;
        f139 = (f139 >= `INH(p234)) ? `INH(p234) : f139;
        f139 = (f139 > p235) ? p235 : f139;
        f140 = 4095;
        f140 = (f140 > p16) ? p16 : f140;
        f140 = (f140 >= `INH(p237)) ? `INH(p237) : f140;
        f141 = 4095;
        f141 = (f141 > p236) ? p236 : f141;
        f141 = (f141 >= `INH(p238)) ? `INH(p238) : f141;
        f142 = 4095;
        f142 = (f142 >= `INH(p16)) ? `INH(p16) : f142;
        f142 = (f142 >= `INH(p237)) ? `INH(p237) : f142;
        f142 = (f142 > p238) ? p238 : f142;
        f143 = 4095;
        f143 = (f143 >= `INH(p236)) ? `INH(p236) : f143;
        f143 = (f143 >= `INH(p238)) ? `INH(p238) : f143;
        f143 = (f143 > p239) ? p239 : f143;
        f144 = 4095;
        f144 = (f144 >= `INH(p5)) ? `INH(p5) : f144;
        f144 = (f144 > p233) ? p233 : f144;
        f144 = (f144 > p237) ? p237 : f144;
        f145 = 4095;
        f145 = (f145 > p219) ? p219 : f145;
        f145 = (f145 >= `INH(p235)) ? `INH(p235) : f145;
        f145 = (f145 >= `INH(p239)) ? `INH(p239) : f145;
        f146 = 4095;
        f146 = (f146 > p220) ? p220 : f146;
        f146 = (f146 >= `INH(p240)) ? `INH(p240) : f146;
        f147 = 4095;
        f147 = (f147 > p17) ? p17 : f147;
        f147 = (f147 >= `INH(p221)) ? `INH(p221) : f147;
        f148 = 4095;
        f148 = (f148 >= `INH(p17)) ? `INH(p17) : f148;
        f148 = (f148 >= `INH(p221)) ? `INH(p221) : f148;
        f148 = (f148 > p240) ? p240 : f148;
        f149 = 4095;
        f149 = (f149 > p6) ? p6 : f149;
        f149 = (f149 >= `INH(p220)) ? `INH(p220) : f149;
        f149 = (f149 >= `INH(p240)) ? `INH(p240) : f149;
        f150 = 4095;
        f150 = (f150 > p242) ? p242 : f150;
        f150 = (f150 >= `INH(p244)) ? `INH(p244) : f150;
        f151 = 4095;
        f151 = (f151 >= `INH(p241)) ? `INH(p241) : f151;
        f151 = (f151 >= `INH(p242)) ? `INH(p242) : f151;
        f151 = (f151 >= `INH(p244)) ? `INH(p244) : f151;
        f151 = (f151 > p245) ? p245 : f151;
        f152 = 4095;
        f152 = (f152 > p14) ? p14 : f152;
        f152 = (f152 >= `INH(p247)) ? `INH(p247) : f152;
        f153 = 4095;
        f153 = (f153 > p246) ? p246 : f153;
        f153 = (f153 >= `INH(p248)) ? `INH(p248) : f153;
        f154 = 4095;
        f154 = (f154 >= `INH(p14)) ? `INH(p14) : f154;
        f154 = (f154 >= `INH(p247)) ? `INH(p247) : f154;
        f154 = (f154 > p248) ? p248 : f154;
        f155 = 4095;
        f155 = (f155 >= `INH(p246)) ? `INH(p246) : f155;
        f155 = (f155 >= `INH(p248)) ? `INH(p248) : f155;
        f155 = (f155 > p249) ? p249 : f155;
        f156 = 4095;
        f156 = (f156 > p17) ? p17 : f156;
        f156 = (f156 >= `INH(p251)) ? `INH(p251) : f156;
        f157 = 4095;
        f157 = (f157 > p250) ? p250 : f157;
        f157 = (f157 >= `INH(p252)) ? `INH(p252) : f157;
        f158 = 4095;
        f158 = (f158 >= `INH(p17)) ? `INH(p17) : f158;
        f158 = (f158 >= `INH(p251)) ? `INH(p251) : f158;
        f158 = (f158 > p252) ? p252 : f158;
        f159 = 4095;
        f159 = (f159 >= `INH(p250)) ? `INH(p250) : f159;
        f159 = (f159 >= `INH(p252)) ? `INH(p252) : f159;
        f159 = (f159 > p253) ? p253 : f159;
        f160 = 4095;
        f160 = (f160 >= `INH(p6)) ? `INH(p6) : f160;
        f160 = (f160 > p247) ? p247 : f160;
        f160 = (f160 > p251) ? p251 : f160;
        f161 = 4095;
        f161 = (f161 > p244) ? p244 : f161;
        f161 = (f161 >= `INH(p249)) ? `INH(p249) : f161;
        f161 = (f161 >= `INH(p253)) ? `INH(p253) : f161;
        f162 = 4095;
        f162 = (f162 > p243) ? p243 : f162;
        f162 = (f162 >= `INH(p254)) ? `INH(p254) : f162;
        f163 = 4095;
        f163 = (f163 > p18) ? p18 : f163;
        f163 = (f163 >= `INH(p245)) ? `INH(p245) : f163;
        f164 = 4095;
        f164 = (f164 >= `INH(p18)) ? `INH(p18) : f164;
        f164 = (f164 >= `INH(p245)) ? `INH(p245) : f164;
        f164 = (f164 > p254) ? p254 : f164;
        f165 = 4095;
        f165 = (f165 > p7) ? p7 : f165;
        f165 = (f165 >= `INH(p243)) ? `INH(p243) : f165;
        f165 = (f165 >= `INH(p254)) ? `INH(p254) : f165;
        f166 = 4095;
        f166 = (f166 >= `INH(p256)) ? `INH(p256) : f166;
        f166 = (f166 >= `INH(p257)) ? `INH(p257) : f166;
        f166 = (f166 > p261) ? p261 : f166;
        f167 = 4095;
        f167 = (f167 > p255) ? p255 : f167;
        f167 = (f167 >= `INH(p261)) ? `INH(p261) : f167;
        f168 = 4095;
        f168 = (f168 > p259) ? p259 : f168;
        f168 = (f168 >= `INH(p261)) ? `INH(p261) : f168;
        f169 = 4095;
        f169 = (f169 >= p256/2) ? p256/2 : f169;
        f169 = (f169 >= `INH(p260)) ? `INH(p260) : f169;
        f170 = 4095;
        f170 = (f170 >= `INH(p260)) ? `INH(p260) : f170;
        f170 = (f170 > p263) ? p263 : f170;
        f171 = 4095;
        f171 = (f171 > p256) ? p256 : f171;
        f171 = (f171 >= `INH(p263)) ? `INH(p263) : f171;
        f171 = (f171 > p265) ? p265 : f171;
        f172 = 4095;
        f172 = (f172 >= `INH(p263)) ? `INH(p263) : f172;
        f172 = (f172 > p266) ? p266 : f172;
        f173 = 4095;
        f173 = (f173 > p255) ? p255 : f173;
        f173 = (f173 >= `INH(p265)) ? `INH(p265) : f173;
        f173 = (f173 >= `INH(p266)) ? `INH(p266) : f173;
        f174 = 4095;
        f174 = (f174 > p255) ? p255 : f174;
        f174 = (f174 >= `INH(p264)) ? `INH(p264) : f174;
        f174 = (f174 >= `INH(p266)) ? `INH(p266) : f174;
        f175 = 4095;
        f175 = (f175 >= `INH(p266)) ? `INH(p266) : f175;
        f175 = (f175 > p268) ? p268 : f175;
        f176 = 4095;
        f176 = (f176 > p262) ? p262 : f176;
        f176 = (f176 >= `INH(p268)) ? `INH(p268) : f176;
        f177 = 4095;
        f177 = (f177 >= `INH(p268)) ? `INH(p268) : f177;
        f177 = (f177 > p269) ? p269 : f177;
        f178 = 4095;
        f178 = (f178 > p267) ? p267 : f178;
        f178 = (f178 >= `INH(p269)) ? `INH(p269) : f178;
        f179 = 4095;
        f179 = (f179 > p257) ? p257 : f179;
        f179 = (f179 > p264) ? p264 : f179;
        f179 = (f179 >= `INH(p265)) ? `INH(p265) : f179;
        f179 = (f179 >= `INH(p269)) ? `INH(p269) : f179;
        f180 = 4095;
        f180 = (f180 > p257) ? p257 : f180;
        f180 = (f180 >= `INH(p264)) ? `INH(p264) : f180;
        f180 = (f180 >= `INH(p269)) ? `INH(p269) : f180;
        f181 = 4095;
        f181 = (f181 > p25) ? p25 : f181;
        f181 = (f181 >= `INH(p271)) ? `INH(p271) : f181;
        f182 = 4095;
        f182 = (f182 > p270) ? p270 : f182;
        f182 = (f182 >= `INH(p272)) ? `INH(p272) : f182;
        f183 = 4095;
        f183 = (f183 >= `INH(p25)) ? `INH(p25) : f183;
        f183 = (f183 >= `INH(p271)) ? `INH(p271) : f183;
        f183 = (f183 > p272) ? p272 : f183;
        f184 = 4095;
        f184 = (f184 >= `INH(p270)) ? `INH(p270) : f184;
        f184 = (f184 >= `INH(p272)) ? `INH(p272) : f184;
        f184 = (f184 > p273) ? p273 : f184;
        f185 = 4095;
        f185 = (f185 > p26) ? p26 : f185;
        f185 = (f185 >= `INH(p275)) ? `INH(p275) : f185;
        f186 = 4095;
        f186 = (f186 > p274) ? p274 : f186;
        f186 = (f186 >= `INH(p276)) ? `INH(p276) : f186;
        f187 = 4095;
        f187 = (f187 >= `INH(p26)) ? `INH(p26) : f187;
        f187 = (f187 >= `INH(p275)) ? `INH(p275) : f187;
        f187 = (f187 > p276) ? p276 : f187;
        f188 = 4095;
        f188 = (f188 >= `INH(p274)) ? `INH(p274) : f188;
        f188 = (f188 >= `INH(p276)) ? `INH(p276) : f188;
        f188 = (f188 > p277) ? p277 : f188;
        f189 = 4095;
        f189 = (f189 >= `INH(p19)) ? `INH(p19) : f189;
        f189 = (f189 > p271) ? p271 : f189;
        f189 = (f189 > p275) ? p275 : f189;
        f190 = 4095;
        f190 = (f190 > p257) ? p257 : f190;
        f190 = (f190 >= `INH(p273)) ? `INH(p273) : f190;
        f190 = (f190 >= `INH(p277)) ? `INH(p277) : f190;
        f191 = 4095;
        f191 = (f191 > p258) ? p258 : f191;
        f191 = (f191 >= `INH(p278)) ? `INH(p278) : f191;
        f192 = 4095;
        f192 = (f192 > p27) ? p27 : f192;
        f192 = (f192 >= `INH(p259)) ? `INH(p259) : f192;
        f193 = 4095;
        f193 = (f193 >= `INH(p27)) ? `INH(p27) : f193;
        f193 = (f193 >= `INH(p259)) ? `INH(p259) : f193;
        f193 = (f193 > p278) ? p278 : f193;
        f194 = 4095;
        f194 = (f194 > p20) ? p20 : f194;
        f194 = (f194 >= `INH(p258)) ? `INH(p258) : f194;
        f194 = (f194 >= `INH(p278)) ? `INH(p278) : f194;
        f195 = 4095;
        f195 = (f195 >= `INH(p280)) ? `INH(p280) : f195;
        f195 = (f195 >= `INH(p281)) ? `INH(p281) : f195;
        f195 = (f195 > p285) ? p285 : f195;
        f196 = 4095;
        f196 = (f196 > p279) ? p279 : f196;
        f196 = (f196 >= `INH(p285)) ? `INH(p285) : f196;
        f197 = 4095;
        f197 = (f197 > p283) ? p283 : f197;
        f197 = (f197 >= `INH(p285)) ? `INH(p285) : f197;
        f198 = 4095;
        f198 = (f198 >= p280/2) ? p280/2 : f198;
        f198 = (f198 >= `INH(p284)) ? `INH(p284) : f198;
        f199 = 4095;
        f199 = (f199 >= `INH(p284)) ? `INH(p284) : f199;
        f199 = (f199 > p287) ? p287 : f199;
        f200 = 4095;
        f200 = (f200 > p280) ? p280 : f200;
        f200 = (f200 >= `INH(p287)) ? `INH(p287) : f200;
        f200 = (f200 > p289) ? p289 : f200;
        f201 = 4095;
        f201 = (f201 >= `INH(p287)) ? `INH(p287) : f201;
        f201 = (f201 > p290) ? p290 : f201;
        f202 = 4095;
        f202 = (f202 > p279) ? p279 : f202;
        f202 = (f202 >= `INH(p289)) ? `INH(p289) : f202;
        f202 = (f202 >= `INH(p290)) ? `INH(p290) : f202;
        f203 = 4095;
        f203 = (f203 > p279) ? p279 : f203;
        f203 = (f203 >= `INH(p288)) ? `INH(p288) : f203;
        f203 = (f203 >= `INH(p290)) ? `INH(p290) : f203;
        f204 = 4095;
        f204 = (f204 >= `INH(p290)) ? `INH(p290) : f204;
        f204 = (f204 > p292) ? p292 : f204;
        f205 = 4095;
        f205 = (f205 > p286) ? p286 : f205;
        f205 = (f205 >= `INH(p292)) ? `INH(p292) : f205;
        f206 = 4095;
        f206 = (f206 >= `INH(p292)) ? `INH(p292) : f206;
        f206 = (f206 > p293) ? p293 : f206;
        f207 = 4095;
        f207 = (f207 > p291) ? p291 : f207;
        f207 = (f207 >= `INH(p293)) ? `INH(p293) : f207;
        f208 = 4095;
        f208 = (f208 > p281) ? p281 : f208;
        f208 = (f208 > p288) ? p288 : f208;
        f208 = (f208 >= `INH(p289)) ? `INH(p289) : f208;
        f208 = (f208 >= `INH(p293)) ? `INH(p293) : f208;
        f209 = 4095;
        f209 = (f209 > p281) ? p281 : f209;
        f209 = (f209 >= `INH(p288)) ? `INH(p288) : f209;
        f209 = (f209 >= `INH(p293)) ? `INH(p293) : f209;
        f210 = 4095;
        f210 = (f210 > p28) ? p28 : f210;
        f210 = (f210 >= `INH(p295)) ? `INH(p295) : f210;
        f211 = 4095;
        f211 = (f211 > p294) ? p294 : f211;
        f211 = (f211 >= `INH(p296)) ? `INH(p296) : f211;
        f212 = 4095;
        f212 = (f212 >= `INH(p28)) ? `INH(p28) : f212;
        f212 = (f212 >= `INH(p295)) ? `INH(p295) : f212;
        f212 = (f212 > p296) ? p296 : f212;
        f213 = 4095;
        f213 = (f213 >= `INH(p294)) ? `INH(p294) : f213;
        f213 = (f213 >= `INH(p296)) ? `INH(p296) : f213;
        f213 = (f213 > p297) ? p297 : f213;
        f214 = 4095;
        f214 = (f214 > p29) ? p29 : f214;
        f214 = (f214 >= `INH(p299)) ? `INH(p299) : f214;
        f215 = 4095;
        f215 = (f215 > p298) ? p298 : f215;
        f215 = (f215 >= `INH(p300)) ? `INH(p300) : f215;
        f216 = 4095;
        f216 = (f216 >= `INH(p29)) ? `INH(p29) : f216;
        f216 = (f216 >= `INH(p299)) ? `INH(p299) : f216;
        f216 = (f216 > p300) ? p300 : f216;
        f217 = 4095;
        f217 = (f217 >= `INH(p298)) ? `INH(p298) : f217;
        f217 = (f217 >= `INH(p300)) ? `INH(p300) : f217;
        f217 = (f217 > p301) ? p301 : f217;
        f218 = 4095;
        f218 = (f218 >= `INH(p20)) ? `INH(p20) : f218;
        f218 = (f218 > p295) ? p295 : f218;
        f218 = (f218 > p299) ? p299 : f218;
        f219 = 4095;
        f219 = (f219 > p281) ? p281 : f219;
        f219 = (f219 >= `INH(p297)) ? `INH(p297) : f219;
        f219 = (f219 >= `INH(p301)) ? `INH(p301) : f219;
        f220 = 4095;
        f220 = (f220 > p282) ? p282 : f220;
        f220 = (f220 >= `INH(p302)) ? `INH(p302) : f220;
        f221 = 4095;
        f221 = (f221 > p30) ? p30 : f221;
        f221 = (f221 >= `INH(p283)) ? `INH(p283) : f221;
        f222 = 4095;
        f222 = (f222 >= `INH(p30)) ? `INH(p30) : f222;
        f222 = (f222 >= `INH(p283)) ? `INH(p283) : f222;
        f222 = (f222 > p302) ? p302 : f222;
        f223 = 4095;
        f223 = (f223 > p21) ? p21 : f223;
        f223 = (f223 >= `INH(p282)) ? `INH(p282) : f223;
        f223 = (f223 >= `INH(p302)) ? `INH(p302) : f223;
        f224 = 4095;
        f224 = (f224 > p304) ? p304 : f224;
        f224 = (f224 >= `INH(p306)) ? `INH(p306) : f224;
        f225 = 4095;
        f225 = (f225 >= `INH(p303)) ? `INH(p303) : f225;
        f225 = (f225 >= `INH(p304)) ? `INH(p304) : f225;
        f225 = (f225 >= `INH(p306)) ? `INH(p306) : f225;
        f225 = (f225 > p307) ? p307 : f225;
        f226 = 4095;
        f226 = (f226 > p27) ? p27 : f226;
        f226 = (f226 >= `INH(p309)) ? `INH(p309) : f226;
        f227 = 4095;
        f227 = (f227 > p308) ? p308 : f227;
        f227 = (f227 >= `INH(p310)) ? `INH(p310) : f227;
        f228 = 4095;
        f228 = (f228 >= `INH(p27)) ? `INH(p27) : f228;
        f228 = (f228 >= `INH(p309)) ? `INH(p309) : f228;
        f228 = (f228 > p310) ? p310 : f228;
        f229 = 4095;
        f229 = (f229 >= `INH(p308)) ? `INH(p308) : f229;
        f229 = (f229 >= `INH(p310)) ? `INH(p310) : f229;
        f229 = (f229 > p311) ? p311 : f229;
        f230 = 4095;
        f230 = (f230 > p30) ? p30 : f230;
        f230 = (f230 >= `INH(p313)) ? `INH(p313) : f230;
        f231 = 4095;
        f231 = (f231 > p312) ? p312 : f231;
        f231 = (f231 >= `INH(p314)) ? `INH(p314) : f231;
        f232 = 4095;
        f232 = (f232 >= `INH(p30)) ? `INH(p30) : f232;
        f232 = (f232 >= `INH(p313)) ? `INH(p313) : f232;
        f232 = (f232 > p314) ? p314 : f232;
        f233 = 4095;
        f233 = (f233 >= `INH(p312)) ? `INH(p312) : f233;
        f233 = (f233 >= `INH(p314)) ? `INH(p314) : f233;
        f233 = (f233 > p315) ? p315 : f233;
        f234 = 4095;
        f234 = (f234 >= `INH(p21)) ? `INH(p21) : f234;
        f234 = (f234 > p309) ? p309 : f234;
        f234 = (f234 > p313) ? p313 : f234;
        f235 = 4095;
        f235 = (f235 > p306) ? p306 : f235;
        f235 = (f235 >= `INH(p311)) ? `INH(p311) : f235;
        f235 = (f235 >= `INH(p315)) ? `INH(p315) : f235;
        f236 = 4095;
        f236 = (f236 > p305) ? p305 : f236;
        f236 = (f236 >= `INH(p316)) ? `INH(p316) : f236;
        f237 = 4095;
        f237 = (f237 > p31) ? p31 : f237;
        f237 = (f237 >= `INH(p307)) ? `INH(p307) : f237;
        f238 = 4095;
        f238 = (f238 >= `INH(p31)) ? `INH(p31) : f238;
        f238 = (f238 >= `INH(p307)) ? `INH(p307) : f238;
        f238 = (f238 > p316) ? p316 : f238;
        f239 = 4095;
        f239 = (f239 > p22) ? p22 : f239;
        f239 = (f239 >= `INH(p305)) ? `INH(p305) : f239;
        f239 = (f239 >= `INH(p316)) ? `INH(p316) : f239;
        f240 = 4095;
        f240 = (f240 >= `INH(p318)) ? `INH(p318) : f240;
        f240 = (f240 >= `INH(p319)) ? `INH(p319) : f240;
        f240 = (f240 > p323) ? p323 : f240;
        f241 = 4095;
        f241 = (f241 > p317) ? p317 : f241;
        f241 = (f241 >= `INH(p323)) ? `INH(p323) : f241;
        f242 = 4095;
        f242 = (f242 > p321) ? p321 : f242;
        f242 = (f242 >= `INH(p323)) ? `INH(p323) : f242;
        f243 = 4095;
        f243 = (f243 >= p318/2) ? p318/2 : f243;
        f243 = (f243 >= `INH(p322)) ? `INH(p322) : f243;
        f244 = 4095;
        f244 = (f244 >= `INH(p322)) ? `INH(p322) : f244;
        f244 = (f244 > p325) ? p325 : f244;
        f245 = 4095;
        f245 = (f245 > p318) ? p318 : f245;
        f245 = (f245 >= `INH(p325)) ? `INH(p325) : f245;
        f245 = (f245 > p327) ? p327 : f245;
        f246 = 4095;
        f246 = (f246 >= `INH(p325)) ? `INH(p325) : f246;
        f246 = (f246 > p328) ? p328 : f246;
        f247 = 4095;
        f247 = (f247 > p317) ? p317 : f247;
        f247 = (f247 >= `INH(p327)) ? `INH(p327) : f247;
        f247 = (f247 >= `INH(p328)) ? `INH(p328) : f247;
        f248 = 4095;
        f248 = (f248 > p317) ? p317 : f248;
        f248 = (f248 >= `INH(p326)) ? `INH(p326) : f248;
        f248 = (f248 >= `INH(p328)) ? `INH(p328) : f248;
        f249 = 4095;
        f249 = (f249 >= `INH(p328)) ? `INH(p328) : f249;
        f249 = (f249 > p330) ? p330 : f249;
        f250 = 4095;
        f250 = (f250 > p324) ? p324 : f250;
        f250 = (f250 >= `INH(p330)) ? `INH(p330) : f250;
        f251 = 4095;
        f251 = (f251 >= `INH(p330)) ? `INH(p330) : f251;
        f251 = (f251 > p331) ? p331 : f251;
        f252 = 4095;
        f252 = (f252 > p329) ? p329 : f252;
        f252 = (f252 >= `INH(p331)) ? `INH(p331) : f252;
        f253 = 4095;
        f253 = (f253 > p319) ? p319 : f253;
        f253 = (f253 > p326) ? p326 : f253;
        f253 = (f253 >= `INH(p327)) ? `INH(p327) : f253;
        f253 = (f253 >= `INH(p331)) ? `INH(p331) : f253;
        f254 = 4095;
        f254 = (f254 > p319) ? p319 : f254;
        f254 = (f254 >= `INH(p326)) ? `INH(p326) : f254;
        f254 = (f254 >= `INH(p331)) ? `INH(p331) : f254;
        f255 = 4095;
        f255 = (f255 > p32) ? p32 : f255;
        f255 = (f255 >= `INH(p333)) ? `INH(p333) : f255;
        f256 = 4095;
        f256 = (f256 > p332) ? p332 : f256;
        f256 = (f256 >= `INH(p334)) ? `INH(p334) : f256;
        f257 = 4095;
        f257 = (f257 >= `INH(p32)) ? `INH(p32) : f257;
        f257 = (f257 >= `INH(p333)) ? `INH(p333) : f257;
        f257 = (f257 > p334) ? p334 : f257;
        f258 = 4095;
        f258 = (f258 >= `INH(p332)) ? `INH(p332) : f258;
        f258 = (f258 >= `INH(p334)) ? `INH(p334) : f258;
        f258 = (f258 > p335) ? p335 : f258;
        f259 = 4095;
        f259 = (f259 > p33) ? p33 : f259;
        f259 = (f259 >= `INH(p337)) ? `INH(p337) : f259;
        f260 = 4095;
        f260 = (f260 > p336) ? p336 : f260;
        f260 = (f260 >= `INH(p338)) ? `INH(p338) : f260;
        f261 = 4095;
        f261 = (f261 >= `INH(p33)) ? `INH(p33) : f261;
        f261 = (f261 >= `INH(p337)) ? `INH(p337) : f261;
        f261 = (f261 > p338) ? p338 : f261;
        f262 = 4095;
        f262 = (f262 >= `INH(p336)) ? `INH(p336) : f262;
        f262 = (f262 >= `INH(p338)) ? `INH(p338) : f262;
        f262 = (f262 > p339) ? p339 : f262;
        f263 = 4095;
        f263 = (f263 >= `INH(p22)) ? `INH(p22) : f263;
        f263 = (f263 > p333) ? p333 : f263;
        f263 = (f263 > p337) ? p337 : f263;
        f264 = 4095;
        f264 = (f264 > p319) ? p319 : f264;
        f264 = (f264 >= `INH(p335)) ? `INH(p335) : f264;
        f264 = (f264 >= `INH(p339)) ? `INH(p339) : f264;
        f265 = 4095;
        f265 = (f265 > p320) ? p320 : f265;
        f265 = (f265 >= `INH(p340)) ? `INH(p340) : f265;
        f266 = 4095;
        f266 = (f266 > p34) ? p34 : f266;
        f266 = (f266 >= `INH(p321)) ? `INH(p321) : f266;
        f267 = 4095;
        f267 = (f267 >= `INH(p34)) ? `INH(p34) : f267;
        f267 = (f267 >= `INH(p321)) ? `INH(p321) : f267;
        f267 = (f267 > p340) ? p340 : f267;
        f268 = 4095;
        f268 = (f268 > p23) ? p23 : f268;
        f268 = (f268 >= `INH(p320)) ? `INH(p320) : f268;
        f268 = (f268 >= `INH(p340)) ? `INH(p340) : f268;
        f269 = 4095;
        f269 = (f269 > p342) ? p342 : f269;
        f269 = (f269 >= `INH(p344)) ? `INH(p344) : f269;
        f270 = 4095;
        f270 = (f270 >= `INH(p341)) ? `INH(p341) : f270;
        f270 = (f270 >= `INH(p342)) ? `INH(p342) : f270;
        f270 = (f270 >= `INH(p344)) ? `INH(p344) : f270;
        f270 = (f270 > p345) ? p345 : f270;
        f271 = 4095;
        f271 = (f271 > p31) ? p31 : f271;
        f271 = (f271 >= `INH(p347)) ? `INH(p347) : f271;
        f272 = 4095;
        f272 = (f272 > p346) ? p346 : f272;
        f272 = (f272 >= `INH(p348)) ? `INH(p348) : f272;
        f273 = 4095;
        f273 = (f273 >= `INH(p31)) ? `INH(p31) : f273;
        f273 = (f273 >= `INH(p347)) ? `INH(p347) : f273;
        f273 = (f273 > p348) ? p348 : f273;
        f274 = 4095;
        f274 = (f274 >= `INH(p346)) ? `INH(p346) : f274;
        f274 = (f274 >= `INH(p348)) ? `INH(p348) : f274;
        f274 = (f274 > p349) ? p349 : f274;
        f275 = 4095;
        f275 = (f275 > p34) ? p34 : f275;
        f275 = (f275 >= `INH(p351)) ? `INH(p351) : f275;
        f276 = 4095;
        f276 = (f276 > p350) ? p350 : f276;
        f276 = (f276 >= `INH(p352)) ? `INH(p352) : f276;
        f277 = 4095;
        f277 = (f277 >= `INH(p34)) ? `INH(p34) : f277;
        f277 = (f277 >= `INH(p351)) ? `INH(p351) : f277;
        f277 = (f277 > p352) ? p352 : f277;
        f278 = 4095;
        f278 = (f278 >= `INH(p350)) ? `INH(p350) : f278;
        f278 = (f278 >= `INH(p352)) ? `INH(p352) : f278;
        f278 = (f278 > p353) ? p353 : f278;
        f279 = 4095;
        f279 = (f279 >= `INH(p23)) ? `INH(p23) : f279;
        f279 = (f279 > p347) ? p347 : f279;
        f279 = (f279 > p351) ? p351 : f279;
        f280 = 4095;
        f280 = (f280 > p344) ? p344 : f280;
        f280 = (f280 >= `INH(p349)) ? `INH(p349) : f280;
        f280 = (f280 >= `INH(p353)) ? `INH(p353) : f280;
        f281 = 4095;
        f281 = (f281 > p343) ? p343 : f281;
        f281 = (f281 >= `INH(p354)) ? `INH(p354) : f281;
        f282 = 4095;
        f282 = (f282 > p35) ? p35 : f282;
        f282 = (f282 >= `INH(p345)) ? `INH(p345) : f282;
        f283 = 4095;
        f283 = (f283 >= `INH(p35)) ? `INH(p35) : f283;
        f283 = (f283 >= `INH(p345)) ? `INH(p345) : f283;
        f283 = (f283 > p354) ? p354 : f283;
        f284 = 4095;
        f284 = (f284 > p24) ? p24 : f284;
        f284 = (f284 >= `INH(p343)) ? `INH(p343) : f284;
        f284 = (f284 >= `INH(p354)) ? `INH(p354) : f284;
        f285 = 4095;
        f285 = (f285 >= `INH(p356)) ? `INH(p356) : f285;
        f285 = (f285 >= `INH(p357)) ? `INH(p357) : f285;
        f285 = (f285 > p361) ? p361 : f285;
        f286 = 4095;
        f286 = (f286 > p355) ? p355 : f286;
        f286 = (f286 >= `INH(p361)) ? `INH(p361) : f286;
        f287 = 4095;
        f287 = (f287 > p359) ? p359 : f287;
        f287 = (f287 >= `INH(p361)) ? `INH(p361) : f287;
        f288 = 4095;
        f288 = (f288 >= p356/2) ? p356/2 : f288;
        f288 = (f288 >= `INH(p360)) ? `INH(p360) : f288;
        f289 = 4095;
        f289 = (f289 >= `INH(p360)) ? `INH(p360) : f289;
        f289 = (f289 > p363) ? p363 : f289;
        f290 = 4095;
        f290 = (f290 > p356) ? p356 : f290;
        f290 = (f290 >= `INH(p363)) ? `INH(p363) : f290;
        f290 = (f290 > p365) ? p365 : f290;
        f291 = 4095;
        f291 = (f291 >= `INH(p363)) ? `INH(p363) : f291;
        f291 = (f291 > p366) ? p366 : f291;
        f292 = 4095;
        f292 = (f292 > p355) ? p355 : f292;
        f292 = (f292 >= `INH(p365)) ? `INH(p365) : f292;
        f292 = (f292 >= `INH(p366)) ? `INH(p366) : f292;
        f293 = 4095;
        f293 = (f293 > p355) ? p355 : f293;
        f293 = (f293 >= `INH(p364)) ? `INH(p364) : f293;
        f293 = (f293 >= `INH(p366)) ? `INH(p366) : f293;
        f294 = 4095;
        f294 = (f294 >= `INH(p366)) ? `INH(p366) : f294;
        f294 = (f294 > p368) ? p368 : f294;
        f295 = 4095;
        f295 = (f295 > p362) ? p362 : f295;
        f295 = (f295 >= `INH(p368)) ? `INH(p368) : f295;
        f296 = 4095;
        f296 = (f296 >= `INH(p368)) ? `INH(p368) : f296;
        f296 = (f296 > p369) ? p369 : f296;
        f297 = 4095;
        f297 = (f297 > p367) ? p367 : f297;
        f297 = (f297 >= `INH(p369)) ? `INH(p369) : f297;
        f298 = 4095;
        f298 = (f298 > p357) ? p357 : f298;
        f298 = (f298 > p364) ? p364 : f298;
        f298 = (f298 >= `INH(p365)) ? `INH(p365) : f298;
        f298 = (f298 >= `INH(p369)) ? `INH(p369) : f298;
        f299 = 4095;
        f299 = (f299 > p357) ? p357 : f299;
        f299 = (f299 >= `INH(p364)) ? `INH(p364) : f299;
        f299 = (f299 >= `INH(p369)) ? `INH(p369) : f299;
        f300 = 4095;
        f300 = (f300 > p42) ? p42 : f300;
        f300 = (f300 >= `INH(p371)) ? `INH(p371) : f300;
        f301 = 4095;
        f301 = (f301 > p370) ? p370 : f301;
        f301 = (f301 >= `INH(p372)) ? `INH(p372) : f301;
        f302 = 4095;
        f302 = (f302 >= `INH(p42)) ? `INH(p42) : f302;
        f302 = (f302 >= `INH(p371)) ? `INH(p371) : f302;
        f302 = (f302 > p372) ? p372 : f302;
        f303 = 4095;
        f303 = (f303 >= `INH(p370)) ? `INH(p370) : f303;
        f303 = (f303 >= `INH(p372)) ? `INH(p372) : f303;
        f303 = (f303 > p373) ? p373 : f303;
        f304 = 4095;
        f304 = (f304 > p43) ? p43 : f304;
        f304 = (f304 >= `INH(p375)) ? `INH(p375) : f304;
        f305 = 4095;
        f305 = (f305 > p374) ? p374 : f305;
        f305 = (f305 >= `INH(p376)) ? `INH(p376) : f305;
        f306 = 4095;
        f306 = (f306 >= `INH(p43)) ? `INH(p43) : f306;
        f306 = (f306 >= `INH(p375)) ? `INH(p375) : f306;
        f306 = (f306 > p376) ? p376 : f306;
        f307 = 4095;
        f307 = (f307 >= `INH(p374)) ? `INH(p374) : f307;
        f307 = (f307 >= `INH(p376)) ? `INH(p376) : f307;
        f307 = (f307 > p377) ? p377 : f307;
        f308 = 4095;
        f308 = (f308 >= `INH(p36)) ? `INH(p36) : f308;
        f308 = (f308 > p371) ? p371 : f308;
        f308 = (f308 > p375) ? p375 : f308;
        f309 = 4095;
        f309 = (f309 > p357) ? p357 : f309;
        f309 = (f309 >= `INH(p373)) ? `INH(p373) : f309;
        f309 = (f309 >= `INH(p377)) ? `INH(p377) : f309;
        f310 = 4095;
        f310 = (f310 > p358) ? p358 : f310;
        f310 = (f310 >= `INH(p378)) ? `INH(p378) : f310;
        f311 = 4095;
        f311 = (f311 > p44) ? p44 : f311;
        f311 = (f311 >= `INH(p359)) ? `INH(p359) : f311;
        f312 = 4095;
        f312 = (f312 >= `INH(p44)) ? `INH(p44) : f312;
        f312 = (f312 >= `INH(p359)) ? `INH(p359) : f312;
        f312 = (f312 > p378) ? p378 : f312;
        f313 = 4095;
        f313 = (f313 > p37) ? p37 : f313;
        f313 = (f313 >= `INH(p358)) ? `INH(p358) : f313;
        f313 = (f313 >= `INH(p378)) ? `INH(p378) : f313;
        f314 = 4095;
        f314 = (f314 >= `INH(p380)) ? `INH(p380) : f314;
        f314 = (f314 >= `INH(p381)) ? `INH(p381) : f314;
        f314 = (f314 > p385) ? p385 : f314;
        f315 = 4095;
        f315 = (f315 > p379) ? p379 : f315;
        f315 = (f315 >= `INH(p385)) ? `INH(p385) : f315;
        f316 = 4095;
        f316 = (f316 > p383) ? p383 : f316;
        f316 = (f316 >= `INH(p385)) ? `INH(p385) : f316;
        f317 = 4095;
        f317 = (f317 >= p380/2) ? p380/2 : f317;
        f317 = (f317 >= `INH(p384)) ? `INH(p384) : f317;
        f318 = 4095;
        f318 = (f318 >= `INH(p384)) ? `INH(p384) : f318;
        f318 = (f318 > p387) ? p387 : f318;
        f319 = 4095;
        f319 = (f319 > p380) ? p380 : f319;
        f319 = (f319 >= `INH(p387)) ? `INH(p387) : f319;
        f319 = (f319 > p389) ? p389 : f319;
        f320 = 4095;
        f320 = (f320 >= `INH(p387)) ? `INH(p387) : f320;
        f320 = (f320 > p390) ? p390 : f320;
        f321 = 4095;
        f321 = (f321 > p379) ? p379 : f321;
        f321 = (f321 >= `INH(p389)) ? `INH(p389) : f321;
        f321 = (f321 >= `INH(p390)) ? `INH(p390) : f321;
        f322 = 4095;
        f322 = (f322 > p379) ? p379 : f322;
        f322 = (f322 >= `INH(p388)) ? `INH(p388) : f322;
        f322 = (f322 >= `INH(p390)) ? `INH(p390) : f322;
        f323 = 4095;
        f323 = (f323 >= `INH(p390)) ? `INH(p390) : f323;
        f323 = (f323 > p392) ? p392 : f323;
        f324 = 4095;
        f324 = (f324 > p386) ? p386 : f324;
        f324 = (f324 >= `INH(p392)) ? `INH(p392) : f324;
        f325 = 4095;
        f325 = (f325 >= `INH(p392)) ? `INH(p392) : f325;
        f325 = (f325 > p393) ? p393 : f325;
        f326 = 4095;
        f326 = (f326 > p391) ? p391 : f326;
        f326 = (f326 >= `INH(p393)) ? `INH(p393) : f326;
        f327 = 4095;
        f327 = (f327 > p381) ? p381 : f327;
        f327 = (f327 > p388) ? p388 : f327;
        f327 = (f327 >= `INH(p389)) ? `INH(p389) : f327;
        f327 = (f327 >= `INH(p393)) ? `INH(p393) : f327;
        f328 = 4095;
        f328 = (f328 > p381) ? p381 : f328;
        f328 = (f328 >= `INH(p388)) ? `INH(p388) : f328;
        f328 = (f328 >= `INH(p393)) ? `INH(p393) : f328;
        f329 = 4095;
        f329 = (f329 > p45) ? p45 : f329;
        f329 = (f329 >= `INH(p395)) ? `INH(p395) : f329;
        f330 = 4095;
        f330 = (f330 > p394) ? p394 : f330;
        f330 = (f330 >= `INH(p396)) ? `INH(p396) : f330;
        f331 = 4095;
        f331 = (f331 >= `INH(p45)) ? `INH(p45) : f331;
        f331 = (f331 >= `INH(p395)) ? `INH(p395) : f331;
        f331 = (f331 > p396) ? p396 : f331;
        f332 = 4095;
        f332 = (f332 >= `INH(p394)) ? `INH(p394) : f332;
        f332 = (f332 >= `INH(p396)) ? `INH(p396) : f332;
        f332 = (f332 > p397) ? p397 : f332;
        f333 = 4095;
        f333 = (f333 > p46) ? p46 : f333;
        f333 = (f333 >= `INH(p399)) ? `INH(p399) : f333;
        f334 = 4095;
        f334 = (f334 > p398) ? p398 : f334;
        f334 = (f334 >= `INH(p400)) ? `INH(p400) : f334;
        f335 = 4095;
        f335 = (f335 >= `INH(p46)) ? `INH(p46) : f335;
        f335 = (f335 >= `INH(p399)) ? `INH(p399) : f335;
        f335 = (f335 > p400) ? p400 : f335;
        f336 = 4095;
        f336 = (f336 >= `INH(p398)) ? `INH(p398) : f336;
        f336 = (f336 >= `INH(p400)) ? `INH(p400) : f336;
        f336 = (f336 > p401) ? p401 : f336;
        f337 = 4095;
        f337 = (f337 >= `INH(p37)) ? `INH(p37) : f337;
        f337 = (f337 > p395) ? p395 : f337;
        f337 = (f337 > p399) ? p399 : f337;
        f338 = 4095;
        f338 = (f338 > p381) ? p381 : f338;
        f338 = (f338 >= `INH(p397)) ? `INH(p397) : f338;
        f338 = (f338 >= `INH(p401)) ? `INH(p401) : f338;
        f339 = 4095;
        f339 = (f339 > p382) ? p382 : f339;
        f339 = (f339 >= `INH(p402)) ? `INH(p402) : f339;
        f340 = 4095;
        f340 = (f340 > p47) ? p47 : f340;
        f340 = (f340 >= `INH(p383)) ? `INH(p383) : f340;
        f341 = 4095;
        f341 = (f341 >= `INH(p47)) ? `INH(p47) : f341;
        f341 = (f341 >= `INH(p383)) ? `INH(p383) : f341;
        f341 = (f341 > p402) ? p402 : f341;
        f342 = 4095;
        f342 = (f342 > p38) ? p38 : f342;
        f342 = (f342 >= `INH(p382)) ? `INH(p382) : f342;
        f342 = (f342 >= `INH(p402)) ? `INH(p402) : f342;
        f343 = 4095;
        f343 = (f343 > p404) ? p404 : f343;
        f343 = (f343 >= `INH(p406)) ? `INH(p406) : f343;
        f344 = 4095;
        f344 = (f344 >= `INH(p403)) ? `INH(p403) : f344;
        f344 = (f344 >= `INH(p404)) ? `INH(p404) : f344;
        f344 = (f344 >= `INH(p406)) ? `INH(p406) : f344;
        f344 = (f344 > p407) ? p407 : f344;
        f345 = 4095;
        f345 = (f345 > p44) ? p44 : f345;
        f345 = (f345 >= `INH(p409)) ? `INH(p409) : f345;
        f346 = 4095;
        f346 = (f346 > p408) ? p408 : f346;
        f346 = (f346 >= `INH(p410)) ? `INH(p410) : f346;
        f347 = 4095;
        f347 = (f347 >= `INH(p44)) ? `INH(p44) : f347;
        f347 = (f347 >= `INH(p409)) ? `INH(p409) : f347;
        f347 = (f347 > p410) ? p410 : f347;
        f348 = 4095;
        f348 = (f348 >= `INH(p408)) ? `INH(p408) : f348;
        f348 = (f348 >= `INH(p410)) ? `INH(p410) : f348;
        f348 = (f348 > p411) ? p411 : f348;
        f349 = 4095;
        f349 = (f349 > p47) ? p47 : f349;
        f349 = (f349 >= `INH(p413)) ? `INH(p413) : f349;
        f350 = 4095;
        f350 = (f350 > p412) ? p412 : f350;
        f350 = (f350 >= `INH(p414)) ? `INH(p414) : f350;
        f351 = 4095;
        f351 = (f351 >= `INH(p47)) ? `INH(p47) : f351;
        f351 = (f351 >= `INH(p413)) ? `INH(p413) : f351;
        f351 = (f351 > p414) ? p414 : f351;
        f352 = 4095;
        f352 = (f352 >= `INH(p412)) ? `INH(p412) : f352;
        f352 = (f352 >= `INH(p414)) ? `INH(p414) : f352;
        f352 = (f352 > p415) ? p415 : f352;
        f353 = 4095;
        f353 = (f353 >= `INH(p38)) ? `INH(p38) : f353;
        f353 = (f353 > p409) ? p409 : f353;
        f353 = (f353 > p413) ? p413 : f353;
        f354 = 4095;
        f354 = (f354 > p406) ? p406 : f354;
        f354 = (f354 >= `INH(p411)) ? `INH(p411) : f354;
        f354 = (f354 >= `INH(p415)) ? `INH(p415) : f354;
        f355 = 4095;
        f355 = (f355 > p405) ? p405 : f355;
        f355 = (f355 >= `INH(p416)) ? `INH(p416) : f355;
        f356 = 4095;
        f356 = (f356 > p48) ? p48 : f356;
        f356 = (f356 >= `INH(p407)) ? `INH(p407) : f356;
        f357 = 4095;
        f357 = (f357 >= `INH(p48)) ? `INH(p48) : f357;
        f357 = (f357 >= `INH(p407)) ? `INH(p407) : f357;
        f357 = (f357 > p416) ? p416 : f357;
        f358 = 4095;
        f358 = (f358 > p39) ? p39 : f358;
        f358 = (f358 >= `INH(p405)) ? `INH(p405) : f358;
        f358 = (f358 >= `INH(p416)) ? `INH(p416) : f358;
        f359 = 4095;
        f359 = (f359 >= `INH(p418)) ? `INH(p418) : f359;
        f359 = (f359 >= `INH(p419)) ? `INH(p419) : f359;
        f359 = (f359 > p423) ? p423 : f359;
        f360 = 4095;
        f360 = (f360 > p417) ? p417 : f360;
        f360 = (f360 >= `INH(p423)) ? `INH(p423) : f360;
        f361 = 4095;
        f361 = (f361 > p421) ? p421 : f361;
        f361 = (f361 >= `INH(p423)) ? `INH(p423) : f361;
        f362 = 4095;
        f362 = (f362 >= p418/2) ? p418/2 : f362;
        f362 = (f362 >= `INH(p422)) ? `INH(p422) : f362;
        f363 = 4095;
        f363 = (f363 >= `INH(p422)) ? `INH(p422) : f363;
        f363 = (f363 > p425) ? p425 : f363;
        f364 = 4095;
        f364 = (f364 > p418) ? p418 : f364;
        f364 = (f364 >= `INH(p425)) ? `INH(p425) : f364;
        f364 = (f364 > p427) ? p427 : f364;
        f365 = 4095;
        f365 = (f365 >= `INH(p425)) ? `INH(p425) : f365;
        f365 = (f365 > p428) ? p428 : f365;
        f366 = 4095;
        f366 = (f366 > p417) ? p417 : f366;
        f366 = (f366 >= `INH(p427)) ? `INH(p427) : f366;
        f366 = (f366 >= `INH(p428)) ? `INH(p428) : f366;
        f367 = 4095;
        f367 = (f367 > p417) ? p417 : f367;
        f367 = (f367 >= `INH(p426)) ? `INH(p426) : f367;
        f367 = (f367 >= `INH(p428)) ? `INH(p428) : f367;
        f368 = 4095;
        f368 = (f368 >= `INH(p428)) ? `INH(p428) : f368;
        f368 = (f368 > p430) ? p430 : f368;
        f369 = 4095;
        f369 = (f369 > p424) ? p424 : f369;
        f369 = (f369 >= `INH(p430)) ? `INH(p430) : f369;
        f370 = 4095;
        f370 = (f370 >= `INH(p430)) ? `INH(p430) : f370;
        f370 = (f370 > p431) ? p431 : f370;
        f371 = 4095;
        f371 = (f371 > p429) ? p429 : f371;
        f371 = (f371 >= `INH(p431)) ? `INH(p431) : f371;
        f372 = 4095;
        f372 = (f372 > p419) ? p419 : f372;
        f372 = (f372 > p426) ? p426 : f372;
        f372 = (f372 >= `INH(p427)) ? `INH(p427) : f372;
        f372 = (f372 >= `INH(p431)) ? `INH(p431) : f372;
        f373 = 4095;
        f373 = (f373 > p419) ? p419 : f373;
        f373 = (f373 >= `INH(p426)) ? `INH(p426) : f373;
        f373 = (f373 >= `INH(p431)) ? `INH(p431) : f373;
        f374 = 4095;
        f374 = (f374 > p49) ? p49 : f374;
        f374 = (f374 >= `INH(p433)) ? `INH(p433) : f374;
        f375 = 4095;
        f375 = (f375 > p432) ? p432 : f375;
        f375 = (f375 >= `INH(p434)) ? `INH(p434) : f375;
        f376 = 4095;
        f376 = (f376 >= `INH(p49)) ? `INH(p49) : f376;
        f376 = (f376 >= `INH(p433)) ? `INH(p433) : f376;
        f376 = (f376 > p434) ? p434 : f376;
        f377 = 4095;
        f377 = (f377 >= `INH(p432)) ? `INH(p432) : f377;
        f377 = (f377 >= `INH(p434)) ? `INH(p434) : f377;
        f377 = (f377 > p435) ? p435 : f377;
        f378 = 4095;
        f378 = (f378 > p50) ? p50 : f378;
        f378 = (f378 >= `INH(p437)) ? `INH(p437) : f378;
        f379 = 4095;
        f379 = (f379 > p436) ? p436 : f379;
        f379 = (f379 >= `INH(p438)) ? `INH(p438) : f379;
        f380 = 4095;
        f380 = (f380 >= `INH(p50)) ? `INH(p50) : f380;
        f380 = (f380 >= `INH(p437)) ? `INH(p437) : f380;
        f380 = (f380 > p438) ? p438 : f380;
        f381 = 4095;
        f381 = (f381 >= `INH(p436)) ? `INH(p436) : f381;
        f381 = (f381 >= `INH(p438)) ? `INH(p438) : f381;
        f381 = (f381 > p439) ? p439 : f381;
        f382 = 4095;
        f382 = (f382 >= `INH(p39)) ? `INH(p39) : f382;
        f382 = (f382 > p433) ? p433 : f382;
        f382 = (f382 > p437) ? p437 : f382;
        f383 = 4095;
        f383 = (f383 > p419) ? p419 : f383;
        f383 = (f383 >= `INH(p435)) ? `INH(p435) : f383;
        f383 = (f383 >= `INH(p439)) ? `INH(p439) : f383;
        f384 = 4095;
        f384 = (f384 > p420) ? p420 : f384;
        f384 = (f384 >= `INH(p440)) ? `INH(p440) : f384;
        f385 = 4095;
        f385 = (f385 > p51) ? p51 : f385;
        f385 = (f385 >= `INH(p421)) ? `INH(p421) : f385;
        f386 = 4095;
        f386 = (f386 >= `INH(p51)) ? `INH(p51) : f386;
        f386 = (f386 >= `INH(p421)) ? `INH(p421) : f386;
        f386 = (f386 > p440) ? p440 : f386;
        f387 = 4095;
        f387 = (f387 > p40) ? p40 : f387;
        f387 = (f387 >= `INH(p420)) ? `INH(p420) : f387;
        f387 = (f387 >= `INH(p440)) ? `INH(p440) : f387;
        f388 = 4095;
        f388 = (f388 > p442) ? p442 : f388;
        f388 = (f388 >= `INH(p444)) ? `INH(p444) : f388;
        f389 = 4095;
        f389 = (f389 >= `INH(p441)) ? `INH(p441) : f389;
        f389 = (f389 >= `INH(p442)) ? `INH(p442) : f389;
        f389 = (f389 >= `INH(p444)) ? `INH(p444) : f389;
        f389 = (f389 > p445) ? p445 : f389;
        f390 = 4095;
        f390 = (f390 > p48) ? p48 : f390;
        f390 = (f390 >= `INH(p447)) ? `INH(p447) : f390;
        f391 = 4095;
        f391 = (f391 > p446) ? p446 : f391;
        f391 = (f391 >= `INH(p448)) ? `INH(p448) : f391;
        f392 = 4095;
        f392 = (f392 >= `INH(p48)) ? `INH(p48) : f392;
        f392 = (f392 >= `INH(p447)) ? `INH(p447) : f392;
        f392 = (f392 > p448) ? p448 : f392;
        f393 = 4095;
        f393 = (f393 >= `INH(p446)) ? `INH(p446) : f393;
        f393 = (f393 >= `INH(p448)) ? `INH(p448) : f393;
        f393 = (f393 > p449) ? p449 : f393;
        f394 = 4095;
        f394 = (f394 > p51) ? p51 : f394;
        f394 = (f394 >= `INH(p451)) ? `INH(p451) : f394;
        f395 = 4095;
        f395 = (f395 > p450) ? p450 : f395;
        f395 = (f395 >= `INH(p452)) ? `INH(p452) : f395;
        f396 = 4095;
        f396 = (f396 >= `INH(p51)) ? `INH(p51) : f396;
        f396 = (f396 >= `INH(p451)) ? `INH(p451) : f396;
        f396 = (f396 > p452) ? p452 : f396;
        f397 = 4095;
        f397 = (f397 >= `INH(p450)) ? `INH(p450) : f397;
        f397 = (f397 >= `INH(p452)) ? `INH(p452) : f397;
        f397 = (f397 > p453) ? p453 : f397;
        f398 = 4095;
        f398 = (f398 >= `INH(p40)) ? `INH(p40) : f398;
        f398 = (f398 > p447) ? p447 : f398;
        f398 = (f398 > p451) ? p451 : f398;
        f399 = 4095;
        f399 = (f399 > p444) ? p444 : f399;
        f399 = (f399 >= `INH(p449)) ? `INH(p449) : f399;
        f399 = (f399 >= `INH(p453)) ? `INH(p453) : f399;
        f400 = 4095;
        f400 = (f400 > p443) ? p443 : f400;
        f400 = (f400 >= `INH(p454)) ? `INH(p454) : f400;
        f401 = 4095;
        f401 = (f401 > p52) ? p52 : f401;
        f401 = (f401 >= `INH(p445)) ? `INH(p445) : f401;
        f402 = 4095;
        f402 = (f402 >= `INH(p52)) ? `INH(p52) : f402;
        f402 = (f402 >= `INH(p445)) ? `INH(p445) : f402;
        f402 = (f402 > p454) ? p454 : f402;
        f403 = 4095;
        f403 = (f403 > p41) ? p41 : f403;
        f403 = (f403 >= `INH(p443)) ? `INH(p443) : f403;
        f403 = (f403 >= `INH(p454)) ? `INH(p454) : f403;
        f404 = 4095;
        f404 = (f404 >= `INH(p456)) ? `INH(p456) : f404;
        f404 = (f404 >= `INH(p457)) ? `INH(p457) : f404;
        f404 = (f404 > p461) ? p461 : f404;
        f405 = 4095;
        f405 = (f405 > p455) ? p455 : f405;
        f405 = (f405 >= `INH(p461)) ? `INH(p461) : f405;
        f406 = 4095;
        f406 = (f406 > p459) ? p459 : f406;
        f406 = (f406 >= `INH(p461)) ? `INH(p461) : f406;
        f407 = 4095;
        f407 = (f407 >= p456/2) ? p456/2 : f407;
        f407 = (f407 >= `INH(p460)) ? `INH(p460) : f407;
        f408 = 4095;
        f408 = (f408 >= `INH(p460)) ? `INH(p460) : f408;
        f408 = (f408 > p463) ? p463 : f408;
        f409 = 4095;
        f409 = (f409 > p456) ? p456 : f409;
        f409 = (f409 >= `INH(p463)) ? `INH(p463) : f409;
        f409 = (f409 > p465) ? p465 : f409;
        f410 = 4095;
        f410 = (f410 >= `INH(p463)) ? `INH(p463) : f410;
        f410 = (f410 > p466) ? p466 : f410;
        f411 = 4095;
        f411 = (f411 > p455) ? p455 : f411;
        f411 = (f411 >= `INH(p465)) ? `INH(p465) : f411;
        f411 = (f411 >= `INH(p466)) ? `INH(p466) : f411;
        f412 = 4095;
        f412 = (f412 > p455) ? p455 : f412;
        f412 = (f412 >= `INH(p464)) ? `INH(p464) : f412;
        f412 = (f412 >= `INH(p466)) ? `INH(p466) : f412;
        f413 = 4095;
        f413 = (f413 >= `INH(p466)) ? `INH(p466) : f413;
        f413 = (f413 > p468) ? p468 : f413;
        f414 = 4095;
        f414 = (f414 > p462) ? p462 : f414;
        f414 = (f414 >= `INH(p468)) ? `INH(p468) : f414;
        f415 = 4095;
        f415 = (f415 >= `INH(p468)) ? `INH(p468) : f415;
        f415 = (f415 > p469) ? p469 : f415;
        f416 = 4095;
        f416 = (f416 > p467) ? p467 : f416;
        f416 = (f416 >= `INH(p469)) ? `INH(p469) : f416;
        f417 = 4095;
        f417 = (f417 > p457) ? p457 : f417;
        f417 = (f417 > p464) ? p464 : f417;
        f417 = (f417 >= `INH(p465)) ? `INH(p465) : f417;
        f417 = (f417 >= `INH(p469)) ? `INH(p469) : f417;
        f418 = 4095;
        f418 = (f418 > p457) ? p457 : f418;
        f418 = (f418 >= `INH(p464)) ? `INH(p464) : f418;
        f418 = (f418 >= `INH(p469)) ? `INH(p469) : f418;
        f419 = 4095;
        f419 = (f419 > p59) ? p59 : f419;
        f419 = (f419 >= `INH(p471)) ? `INH(p471) : f419;
        f420 = 4095;
        f420 = (f420 > p470) ? p470 : f420;
        f420 = (f420 >= `INH(p472)) ? `INH(p472) : f420;
        f421 = 4095;
        f421 = (f421 >= `INH(p59)) ? `INH(p59) : f421;
        f421 = (f421 >= `INH(p471)) ? `INH(p471) : f421;
        f421 = (f421 > p472) ? p472 : f421;
        f422 = 4095;
        f422 = (f422 >= `INH(p470)) ? `INH(p470) : f422;
        f422 = (f422 >= `INH(p472)) ? `INH(p472) : f422;
        f422 = (f422 > p473) ? p473 : f422;
        f423 = 4095;
        f423 = (f423 > p60) ? p60 : f423;
        f423 = (f423 >= `INH(p475)) ? `INH(p475) : f423;
        f424 = 4095;
        f424 = (f424 > p474) ? p474 : f424;
        f424 = (f424 >= `INH(p476)) ? `INH(p476) : f424;
        f425 = 4095;
        f425 = (f425 >= `INH(p60)) ? `INH(p60) : f425;
        f425 = (f425 >= `INH(p475)) ? `INH(p475) : f425;
        f425 = (f425 > p476) ? p476 : f425;
        f426 = 4095;
        f426 = (f426 >= `INH(p474)) ? `INH(p474) : f426;
        f426 = (f426 >= `INH(p476)) ? `INH(p476) : f426;
        f426 = (f426 > p477) ? p477 : f426;
        f427 = 4095;
        f427 = (f427 >= `INH(p53)) ? `INH(p53) : f427;
        f427 = (f427 > p471) ? p471 : f427;
        f427 = (f427 > p475) ? p475 : f427;
        f428 = 4095;
        f428 = (f428 > p457) ? p457 : f428;
        f428 = (f428 >= `INH(p473)) ? `INH(p473) : f428;
        f428 = (f428 >= `INH(p477)) ? `INH(p477) : f428;
        f429 = 4095;
        f429 = (f429 > p458) ? p458 : f429;
        f429 = (f429 >= `INH(p478)) ? `INH(p478) : f429;
        f430 = 4095;
        f430 = (f430 > p61) ? p61 : f430;
        f430 = (f430 >= `INH(p459)) ? `INH(p459) : f430;
        f431 = 4095;
        f431 = (f431 >= `INH(p61)) ? `INH(p61) : f431;
        f431 = (f431 >= `INH(p459)) ? `INH(p459) : f431;
        f431 = (f431 > p478) ? p478 : f431;
        f432 = 4095;
        f432 = (f432 > p54) ? p54 : f432;
        f432 = (f432 >= `INH(p458)) ? `INH(p458) : f432;
        f432 = (f432 >= `INH(p478)) ? `INH(p478) : f432;
        f433 = 4095;
        f433 = (f433 >= `INH(p480)) ? `INH(p480) : f433;
        f433 = (f433 >= `INH(p481)) ? `INH(p481) : f433;
        f433 = (f433 > p485) ? p485 : f433;
        f434 = 4095;
        f434 = (f434 > p479) ? p479 : f434;
        f434 = (f434 >= `INH(p485)) ? `INH(p485) : f434;
        f435 = 4095;
        f435 = (f435 > p483) ? p483 : f435;
        f435 = (f435 >= `INH(p485)) ? `INH(p485) : f435;
        f436 = 4095;
        f436 = (f436 >= p480/2) ? p480/2 : f436;
        f436 = (f436 >= `INH(p484)) ? `INH(p484) : f436;
        f437 = 4095;
        f437 = (f437 >= `INH(p484)) ? `INH(p484) : f437;
        f437 = (f437 > p487) ? p487 : f437;
        f438 = 4095;
        f438 = (f438 > p480) ? p480 : f438;
        f438 = (f438 >= `INH(p487)) ? `INH(p487) : f438;
        f438 = (f438 > p489) ? p489 : f438;
        f439 = 4095;
        f439 = (f439 >= `INH(p487)) ? `INH(p487) : f439;
        f439 = (f439 > p490) ? p490 : f439;
        f440 = 4095;
        f440 = (f440 > p479) ? p479 : f440;
        f440 = (f440 >= `INH(p489)) ? `INH(p489) : f440;
        f440 = (f440 >= `INH(p490)) ? `INH(p490) : f440;
        f441 = 4095;
        f441 = (f441 > p479) ? p479 : f441;
        f441 = (f441 >= `INH(p488)) ? `INH(p488) : f441;
        f441 = (f441 >= `INH(p490)) ? `INH(p490) : f441;
        f442 = 4095;
        f442 = (f442 >= `INH(p490)) ? `INH(p490) : f442;
        f442 = (f442 > p492) ? p492 : f442;
        f443 = 4095;
        f443 = (f443 > p486) ? p486 : f443;
        f443 = (f443 >= `INH(p492)) ? `INH(p492) : f443;
        f444 = 4095;
        f444 = (f444 >= `INH(p492)) ? `INH(p492) : f444;
        f444 = (f444 > p493) ? p493 : f444;
        f445 = 4095;
        f445 = (f445 > p491) ? p491 : f445;
        f445 = (f445 >= `INH(p493)) ? `INH(p493) : f445;
        f446 = 4095;
        f446 = (f446 > p481) ? p481 : f446;
        f446 = (f446 > p488) ? p488 : f446;
        f446 = (f446 >= `INH(p489)) ? `INH(p489) : f446;
        f446 = (f446 >= `INH(p493)) ? `INH(p493) : f446;
        f447 = 4095;
        f447 = (f447 > p481) ? p481 : f447;
        f447 = (f447 >= `INH(p488)) ? `INH(p488) : f447;
        f447 = (f447 >= `INH(p493)) ? `INH(p493) : f447;
        f448 = 4095;
        f448 = (f448 > p62) ? p62 : f448;
        f448 = (f448 >= `INH(p495)) ? `INH(p495) : f448;
        f449 = 4095;
        f449 = (f449 > p494) ? p494 : f449;
        f449 = (f449 >= `INH(p496)) ? `INH(p496) : f449;
        f450 = 4095;
        f450 = (f450 >= `INH(p62)) ? `INH(p62) : f450;
        f450 = (f450 >= `INH(p495)) ? `INH(p495) : f450;
        f450 = (f450 > p496) ? p496 : f450;
        f451 = 4095;
        f451 = (f451 >= `INH(p494)) ? `INH(p494) : f451;
        f451 = (f451 >= `INH(p496)) ? `INH(p496) : f451;
        f451 = (f451 > p497) ? p497 : f451;
        f452 = 4095;
        f452 = (f452 > p63) ? p63 : f452;
        f452 = (f452 >= `INH(p499)) ? `INH(p499) : f452;
        f453 = 4095;
        f453 = (f453 > p498) ? p498 : f453;
        f453 = (f453 >= `INH(p500)) ? `INH(p500) : f453;
        f454 = 4095;
        f454 = (f454 >= `INH(p63)) ? `INH(p63) : f454;
        f454 = (f454 >= `INH(p499)) ? `INH(p499) : f454;
        f454 = (f454 > p500) ? p500 : f454;
        f455 = 4095;
        f455 = (f455 >= `INH(p498)) ? `INH(p498) : f455;
        f455 = (f455 >= `INH(p500)) ? `INH(p500) : f455;
        f455 = (f455 > p501) ? p501 : f455;
        f456 = 4095;
        f456 = (f456 >= `INH(p54)) ? `INH(p54) : f456;
        f456 = (f456 > p495) ? p495 : f456;
        f456 = (f456 > p499) ? p499 : f456;
        f457 = 4095;
        f457 = (f457 > p481) ? p481 : f457;
        f457 = (f457 >= `INH(p497)) ? `INH(p497) : f457;
        f457 = (f457 >= `INH(p501)) ? `INH(p501) : f457;
        f458 = 4095;
        f458 = (f458 > p482) ? p482 : f458;
        f458 = (f458 >= `INH(p502)) ? `INH(p502) : f458;
        f459 = 4095;
        f459 = (f459 > p64) ? p64 : f459;
        f459 = (f459 >= `INH(p483)) ? `INH(p483) : f459;
        f460 = 4095;
        f460 = (f460 >= `INH(p64)) ? `INH(p64) : f460;
        f460 = (f460 >= `INH(p483)) ? `INH(p483) : f460;
        f460 = (f460 > p502) ? p502 : f460;
        f461 = 4095;
        f461 = (f461 > p55) ? p55 : f461;
        f461 = (f461 >= `INH(p482)) ? `INH(p482) : f461;
        f461 = (f461 >= `INH(p502)) ? `INH(p502) : f461;
        f462 = 4095;
        f462 = (f462 > p504) ? p504 : f462;
        f462 = (f462 >= `INH(p506)) ? `INH(p506) : f462;
        f463 = 4095;
        f463 = (f463 >= `INH(p503)) ? `INH(p503) : f463;
        f463 = (f463 >= `INH(p504)) ? `INH(p504) : f463;
        f463 = (f463 >= `INH(p506)) ? `INH(p506) : f463;
        f463 = (f463 > p507) ? p507 : f463;
        f464 = 4095;
        f464 = (f464 > p61) ? p61 : f464;
        f464 = (f464 >= `INH(p509)) ? `INH(p509) : f464;
        f465 = 4095;
        f465 = (f465 > p508) ? p508 : f465;
        f465 = (f465 >= `INH(p510)) ? `INH(p510) : f465;
        f466 = 4095;
        f466 = (f466 >= `INH(p61)) ? `INH(p61) : f466;
        f466 = (f466 >= `INH(p509)) ? `INH(p509) : f466;
        f466 = (f466 > p510) ? p510 : f466;
        f467 = 4095;
        f467 = (f467 >= `INH(p508)) ? `INH(p508) : f467;
        f467 = (f467 >= `INH(p510)) ? `INH(p510) : f467;
        f467 = (f467 > p511) ? p511 : f467;
        f468 = 4095;
        f468 = (f468 > p64) ? p64 : f468;
        f468 = (f468 >= `INH(p513)) ? `INH(p513) : f468;
        f469 = 4095;
        f469 = (f469 > p512) ? p512 : f469;
        f469 = (f469 >= `INH(p514)) ? `INH(p514) : f469;
        f470 = 4095;
        f470 = (f470 >= `INH(p64)) ? `INH(p64) : f470;
        f470 = (f470 >= `INH(p513)) ? `INH(p513) : f470;
        f470 = (f470 > p514) ? p514 : f470;
        f471 = 4095;
        f471 = (f471 >= `INH(p512)) ? `INH(p512) : f471;
        f471 = (f471 >= `INH(p514)) ? `INH(p514) : f471;
        f471 = (f471 > p515) ? p515 : f471;
        f472 = 4095;
        f472 = (f472 >= `INH(p55)) ? `INH(p55) : f472;
        f472 = (f472 > p509) ? p509 : f472;
        f472 = (f472 > p513) ? p513 : f472;
        f473 = 4095;
        f473 = (f473 > p506) ? p506 : f473;
        f473 = (f473 >= `INH(p511)) ? `INH(p511) : f473;
        f473 = (f473 >= `INH(p515)) ? `INH(p515) : f473;
        f474 = 4095;
        f474 = (f474 > p505) ? p505 : f474;
        f474 = (f474 >= `INH(p516)) ? `INH(p516) : f474;
        f475 = 4095;
        f475 = (f475 > p65) ? p65 : f475;
        f475 = (f475 >= `INH(p507)) ? `INH(p507) : f475;
        f476 = 4095;
        f476 = (f476 >= `INH(p65)) ? `INH(p65) : f476;
        f476 = (f476 >= `INH(p507)) ? `INH(p507) : f476;
        f476 = (f476 > p516) ? p516 : f476;
        f477 = 4095;
        f477 = (f477 > p56) ? p56 : f477;
        f477 = (f477 >= `INH(p505)) ? `INH(p505) : f477;
        f477 = (f477 >= `INH(p516)) ? `INH(p516) : f477;
        f478 = 4095;
        f478 = (f478 >= `INH(p518)) ? `INH(p518) : f478;
        f478 = (f478 >= `INH(p519)) ? `INH(p519) : f478;
        f478 = (f478 > p523) ? p523 : f478;
        f479 = 4095;
        f479 = (f479 > p517) ? p517 : f479;
        f479 = (f479 >= `INH(p523)) ? `INH(p523) : f479;
        f480 = 4095;
        f480 = (f480 > p521) ? p521 : f480;
        f480 = (f480 >= `INH(p523)) ? `INH(p523) : f480;
        f481 = 4095;
        f481 = (f481 >= p518/2) ? p518/2 : f481;
        f481 = (f481 >= `INH(p522)) ? `INH(p522) : f481;
        f482 = 4095;
        f482 = (f482 >= `INH(p522)) ? `INH(p522) : f482;
        f482 = (f482 > p525) ? p525 : f482;
        f483 = 4095;
        f483 = (f483 > p518) ? p518 : f483;
        f483 = (f483 >= `INH(p525)) ? `INH(p525) : f483;
        f483 = (f483 > p527) ? p527 : f483;
        f484 = 4095;
        f484 = (f484 >= `INH(p525)) ? `INH(p525) : f484;
        f484 = (f484 > p528) ? p528 : f484;
        f485 = 4095;
        f485 = (f485 > p517) ? p517 : f485;
        f485 = (f485 >= `INH(p527)) ? `INH(p527) : f485;
        f485 = (f485 >= `INH(p528)) ? `INH(p528) : f485;
        f486 = 4095;
        f486 = (f486 > p517) ? p517 : f486;
        f486 = (f486 >= `INH(p526)) ? `INH(p526) : f486;
        f486 = (f486 >= `INH(p528)) ? `INH(p528) : f486;
        f487 = 4095;
        f487 = (f487 >= `INH(p528)) ? `INH(p528) : f487;
        f487 = (f487 > p530) ? p530 : f487;
        f488 = 4095;
        f488 = (f488 > p524) ? p524 : f488;
        f488 = (f488 >= `INH(p530)) ? `INH(p530) : f488;
        f489 = 4095;
        f489 = (f489 >= `INH(p530)) ? `INH(p530) : f489;
        f489 = (f489 > p531) ? p531 : f489;
        f490 = 4095;
        f490 = (f490 > p529) ? p529 : f490;
        f490 = (f490 >= `INH(p531)) ? `INH(p531) : f490;
        f491 = 4095;
        f491 = (f491 > p519) ? p519 : f491;
        f491 = (f491 > p526) ? p526 : f491;
        f491 = (f491 >= `INH(p527)) ? `INH(p527) : f491;
        f491 = (f491 >= `INH(p531)) ? `INH(p531) : f491;
        f492 = 4095;
        f492 = (f492 > p519) ? p519 : f492;
        f492 = (f492 >= `INH(p526)) ? `INH(p526) : f492;
        f492 = (f492 >= `INH(p531)) ? `INH(p531) : f492;
        f493 = 4095;
        f493 = (f493 > p66) ? p66 : f493;
        f493 = (f493 >= `INH(p533)) ? `INH(p533) : f493;
        f494 = 4095;
        f494 = (f494 > p532) ? p532 : f494;
        f494 = (f494 >= `INH(p534)) ? `INH(p534) : f494;
        f495 = 4095;
        f495 = (f495 >= `INH(p66)) ? `INH(p66) : f495;
        f495 = (f495 >= `INH(p533)) ? `INH(p533) : f495;
        f495 = (f495 > p534) ? p534 : f495;
        f496 = 4095;
        f496 = (f496 >= `INH(p532)) ? `INH(p532) : f496;
        f496 = (f496 >= `INH(p534)) ? `INH(p534) : f496;
        f496 = (f496 > p535) ? p535 : f496;
        f497 = 4095;
        f497 = (f497 > p67) ? p67 : f497;
        f497 = (f497 >= `INH(p537)) ? `INH(p537) : f497;
        f498 = 4095;
        f498 = (f498 > p536) ? p536 : f498;
        f498 = (f498 >= `INH(p538)) ? `INH(p538) : f498;
        f499 = 4095;
        f499 = (f499 >= `INH(p67)) ? `INH(p67) : f499;
        f499 = (f499 >= `INH(p537)) ? `INH(p537) : f499;
        f499 = (f499 > p538) ? p538 : f499;
        f500 = 4095;
        f500 = (f500 >= `INH(p536)) ? `INH(p536) : f500;
        f500 = (f500 >= `INH(p538)) ? `INH(p538) : f500;
        f500 = (f500 > p539) ? p539 : f500;
        f501 = 4095;
        f501 = (f501 >= `INH(p56)) ? `INH(p56) : f501;
        f501 = (f501 > p533) ? p533 : f501;
        f501 = (f501 > p537) ? p537 : f501;
        f502 = 4095;
        f502 = (f502 > p519) ? p519 : f502;
        f502 = (f502 >= `INH(p535)) ? `INH(p535) : f502;
        f502 = (f502 >= `INH(p539)) ? `INH(p539) : f502;
        f503 = 4095;
        f503 = (f503 > p520) ? p520 : f503;
        f503 = (f503 >= `INH(p540)) ? `INH(p540) : f503;
        f504 = 4095;
        f504 = (f504 > p68) ? p68 : f504;
        f504 = (f504 >= `INH(p521)) ? `INH(p521) : f504;
        f505 = 4095;
        f505 = (f505 >= `INH(p68)) ? `INH(p68) : f505;
        f505 = (f505 >= `INH(p521)) ? `INH(p521) : f505;
        f505 = (f505 > p540) ? p540 : f505;
        f506 = 4095;
        f506 = (f506 > p57) ? p57 : f506;
        f506 = (f506 >= `INH(p520)) ? `INH(p520) : f506;
        f506 = (f506 >= `INH(p540)) ? `INH(p540) : f506;
        f507 = 4095;
        f507 = (f507 > p542) ? p542 : f507;
        f507 = (f507 >= `INH(p544)) ? `INH(p544) : f507;
        f508 = 4095;
        f508 = (f508 >= `INH(p541)) ? `INH(p541) : f508;
        f508 = (f508 >= `INH(p542)) ? `INH(p542) : f508;
        f508 = (f508 >= `INH(p544)) ? `INH(p544) : f508;
        f508 = (f508 > p545) ? p545 : f508;
        f509 = 4095;
        f509 = (f509 > p65) ? p65 : f509;
        f509 = (f509 >= `INH(p547)) ? `INH(p547) : f509;
        f510 = 4095;
        f510 = (f510 > p546) ? p546 : f510;
        f510 = (f510 >= `INH(p548)) ? `INH(p548) : f510;
        f511 = 4095;
        f511 = (f511 >= `INH(p65)) ? `INH(p65) : f511;
        f511 = (f511 >= `INH(p547)) ? `INH(p547) : f511;
        f511 = (f511 > p548) ? p548 : f511;
        f512 = 4095;
        f512 = (f512 >= `INH(p546)) ? `INH(p546) : f512;
        f512 = (f512 >= `INH(p548)) ? `INH(p548) : f512;
        f512 = (f512 > p549) ? p549 : f512;
        f513 = 4095;
        f513 = (f513 > p68) ? p68 : f513;
        f513 = (f513 >= `INH(p551)) ? `INH(p551) : f513;
        f514 = 4095;
        f514 = (f514 > p550) ? p550 : f514;
        f514 = (f514 >= `INH(p552)) ? `INH(p552) : f514;
        f515 = 4095;
        f515 = (f515 >= `INH(p68)) ? `INH(p68) : f515;
        f515 = (f515 >= `INH(p551)) ? `INH(p551) : f515;
        f515 = (f515 > p552) ? p552 : f515;
        f516 = 4095;
        f516 = (f516 >= `INH(p550)) ? `INH(p550) : f516;
        f516 = (f516 >= `INH(p552)) ? `INH(p552) : f516;
        f516 = (f516 > p553) ? p553 : f516;
        f517 = 4095;
        f517 = (f517 >= `INH(p57)) ? `INH(p57) : f517;
        f517 = (f517 > p547) ? p547 : f517;
        f517 = (f517 > p551) ? p551 : f517;
        f518 = 4095;
        f518 = (f518 > p544) ? p544 : f518;
        f518 = (f518 >= `INH(p549)) ? `INH(p549) : f518;
        f518 = (f518 >= `INH(p553)) ? `INH(p553) : f518;
        f519 = 4095;
        f519 = (f519 > p543) ? p543 : f519;
        f519 = (f519 >= `INH(p554)) ? `INH(p554) : f519;
        f520 = 4095;
        f520 = (f520 > p69) ? p69 : f520;
        f520 = (f520 >= `INH(p545)) ? `INH(p545) : f520;
        f521 = 4095;
        f521 = (f521 >= `INH(p69)) ? `INH(p69) : f521;
        f521 = (f521 >= `INH(p545)) ? `INH(p545) : f521;
        f521 = (f521 > p554) ? p554 : f521;
        f522 = 4095;
        f522 = (f522 > p58) ? p58 : f522;
        f522 = (f522 >= `INH(p543)) ? `INH(p543) : f522;
        f522 = (f522 >= `INH(p554)) ? `INH(p554) : f522;
        f523 = 4095;
        f523 = (f523 >= `INH(p556)) ? `INH(p556) : f523;
        f523 = (f523 >= `INH(p557)) ? `INH(p557) : f523;
        f523 = (f523 > p561) ? p561 : f523;
        f524 = 4095;
        f524 = (f524 > p555) ? p555 : f524;
        f524 = (f524 >= `INH(p561)) ? `INH(p561) : f524;
        f525 = 4095;
        f525 = (f525 > p559) ? p559 : f525;
        f525 = (f525 >= `INH(p561)) ? `INH(p561) : f525;
        f526 = 4095;
        f526 = (f526 >= p556/2) ? p556/2 : f526;
        f526 = (f526 >= `INH(p560)) ? `INH(p560) : f526;
        f527 = 4095;
        f527 = (f527 >= `INH(p560)) ? `INH(p560) : f527;
        f527 = (f527 > p563) ? p563 : f527;
        f528 = 4095;
        f528 = (f528 > p556) ? p556 : f528;
        f528 = (f528 >= `INH(p563)) ? `INH(p563) : f528;
        f528 = (f528 > p565) ? p565 : f528;
        f529 = 4095;
        f529 = (f529 >= `INH(p563)) ? `INH(p563) : f529;
        f529 = (f529 > p566) ? p566 : f529;
        f530 = 4095;
        f530 = (f530 > p555) ? p555 : f530;
        f530 = (f530 >= `INH(p565)) ? `INH(p565) : f530;
        f530 = (f530 >= `INH(p566)) ? `INH(p566) : f530;
        f531 = 4095;
        f531 = (f531 > p555) ? p555 : f531;
        f531 = (f531 >= `INH(p564)) ? `INH(p564) : f531;
        f531 = (f531 >= `INH(p566)) ? `INH(p566) : f531;
        f532 = 4095;
        f532 = (f532 >= `INH(p566)) ? `INH(p566) : f532;
        f532 = (f532 > p568) ? p568 : f532;
        f533 = 4095;
        f533 = (f533 > p562) ? p562 : f533;
        f533 = (f533 >= `INH(p568)) ? `INH(p568) : f533;
        f534 = 4095;
        f534 = (f534 >= `INH(p568)) ? `INH(p568) : f534;
        f534 = (f534 > p569) ? p569 : f534;
        f535 = 4095;
        f535 = (f535 > p567) ? p567 : f535;
        f535 = (f535 >= `INH(p569)) ? `INH(p569) : f535;
        f536 = 4095;
        f536 = (f536 > p557) ? p557 : f536;
        f536 = (f536 > p564) ? p564 : f536;
        f536 = (f536 >= `INH(p565)) ? `INH(p565) : f536;
        f536 = (f536 >= `INH(p569)) ? `INH(p569) : f536;
        f537 = 4095;
        f537 = (f537 > p557) ? p557 : f537;
        f537 = (f537 >= `INH(p564)) ? `INH(p564) : f537;
        f537 = (f537 >= `INH(p569)) ? `INH(p569) : f537;
        f538 = 4095;
        f538 = (f538 > p76) ? p76 : f538;
        f538 = (f538 >= `INH(p571)) ? `INH(p571) : f538;
        f539 = 4095;
        f539 = (f539 > p570) ? p570 : f539;
        f539 = (f539 >= `INH(p572)) ? `INH(p572) : f539;
        f540 = 4095;
        f540 = (f540 >= `INH(p76)) ? `INH(p76) : f540;
        f540 = (f540 >= `INH(p571)) ? `INH(p571) : f540;
        f540 = (f540 > p572) ? p572 : f540;
        f541 = 4095;
        f541 = (f541 >= `INH(p570)) ? `INH(p570) : f541;
        f541 = (f541 >= `INH(p572)) ? `INH(p572) : f541;
        f541 = (f541 > p573) ? p573 : f541;
        f542 = 4095;
        f542 = (f542 > p77) ? p77 : f542;
        f542 = (f542 >= `INH(p575)) ? `INH(p575) : f542;
        f543 = 4095;
        f543 = (f543 > p574) ? p574 : f543;
        f543 = (f543 >= `INH(p576)) ? `INH(p576) : f543;
        f544 = 4095;
        f544 = (f544 >= `INH(p77)) ? `INH(p77) : f544;
        f544 = (f544 >= `INH(p575)) ? `INH(p575) : f544;
        f544 = (f544 > p576) ? p576 : f544;
        f545 = 4095;
        f545 = (f545 >= `INH(p574)) ? `INH(p574) : f545;
        f545 = (f545 >= `INH(p576)) ? `INH(p576) : f545;
        f545 = (f545 > p577) ? p577 : f545;
        f546 = 4095;
        f546 = (f546 >= `INH(p70)) ? `INH(p70) : f546;
        f546 = (f546 > p571) ? p571 : f546;
        f546 = (f546 > p575) ? p575 : f546;
        f547 = 4095;
        f547 = (f547 > p557) ? p557 : f547;
        f547 = (f547 >= `INH(p573)) ? `INH(p573) : f547;
        f547 = (f547 >= `INH(p577)) ? `INH(p577) : f547;
        f548 = 4095;
        f548 = (f548 > p558) ? p558 : f548;
        f548 = (f548 >= `INH(p578)) ? `INH(p578) : f548;
        f549 = 4095;
        f549 = (f549 > p78) ? p78 : f549;
        f549 = (f549 >= `INH(p559)) ? `INH(p559) : f549;
        f550 = 4095;
        f550 = (f550 >= `INH(p78)) ? `INH(p78) : f550;
        f550 = (f550 >= `INH(p559)) ? `INH(p559) : f550;
        f550 = (f550 > p578) ? p578 : f550;
        f551 = 4095;
        f551 = (f551 > p71) ? p71 : f551;
        f551 = (f551 >= `INH(p558)) ? `INH(p558) : f551;
        f551 = (f551 >= `INH(p578)) ? `INH(p578) : f551;
        f552 = 4095;
        f552 = (f552 >= `INH(p580)) ? `INH(p580) : f552;
        f552 = (f552 >= `INH(p581)) ? `INH(p581) : f552;
        f552 = (f552 > p585) ? p585 : f552;
        f553 = 4095;
        f553 = (f553 > p579) ? p579 : f553;
        f553 = (f553 >= `INH(p585)) ? `INH(p585) : f553;
        f554 = 4095;
        f554 = (f554 > p583) ? p583 : f554;
        f554 = (f554 >= `INH(p585)) ? `INH(p585) : f554;
        f555 = 4095;
        f555 = (f555 >= p580/2) ? p580/2 : f555;
        f555 = (f555 >= `INH(p584)) ? `INH(p584) : f555;
        f556 = 4095;
        f556 = (f556 >= `INH(p584)) ? `INH(p584) : f556;
        f556 = (f556 > p587) ? p587 : f556;
        f557 = 4095;
        f557 = (f557 > p580) ? p580 : f557;
        f557 = (f557 >= `INH(p587)) ? `INH(p587) : f557;
        f557 = (f557 > p589) ? p589 : f557;
        f558 = 4095;
        f558 = (f558 >= `INH(p587)) ? `INH(p587) : f558;
        f558 = (f558 > p590) ? p590 : f558;
        f559 = 4095;
        f559 = (f559 > p579) ? p579 : f559;
        f559 = (f559 >= `INH(p589)) ? `INH(p589) : f559;
        f559 = (f559 >= `INH(p590)) ? `INH(p590) : f559;
        f560 = 4095;
        f560 = (f560 > p579) ? p579 : f560;
        f560 = (f560 >= `INH(p588)) ? `INH(p588) : f560;
        f560 = (f560 >= `INH(p590)) ? `INH(p590) : f560;
        f561 = 4095;
        f561 = (f561 >= `INH(p590)) ? `INH(p590) : f561;
        f561 = (f561 > p592) ? p592 : f561;
        f562 = 4095;
        f562 = (f562 > p586) ? p586 : f562;
        f562 = (f562 >= `INH(p592)) ? `INH(p592) : f562;
        f563 = 4095;
        f563 = (f563 >= `INH(p592)) ? `INH(p592) : f563;
        f563 = (f563 > p593) ? p593 : f563;
        f564 = 4095;
        f564 = (f564 > p591) ? p591 : f564;
        f564 = (f564 >= `INH(p593)) ? `INH(p593) : f564;
        f565 = 4095;
        f565 = (f565 > p581) ? p581 : f565;
        f565 = (f565 > p588) ? p588 : f565;
        f565 = (f565 >= `INH(p589)) ? `INH(p589) : f565;
        f565 = (f565 >= `INH(p593)) ? `INH(p593) : f565;
        f566 = 4095;
        f566 = (f566 > p581) ? p581 : f566;
        f566 = (f566 >= `INH(p588)) ? `INH(p588) : f566;
        f566 = (f566 >= `INH(p593)) ? `INH(p593) : f566;
        f567 = 4095;
        f567 = (f567 > p79) ? p79 : f567;
        f567 = (f567 >= `INH(p595)) ? `INH(p595) : f567;
        f568 = 4095;
        f568 = (f568 > p594) ? p594 : f568;
        f568 = (f568 >= `INH(p596)) ? `INH(p596) : f568;
        f569 = 4095;
        f569 = (f569 >= `INH(p79)) ? `INH(p79) : f569;
        f569 = (f569 >= `INH(p595)) ? `INH(p595) : f569;
        f569 = (f569 > p596) ? p596 : f569;
        f570 = 4095;
        f570 = (f570 >= `INH(p594)) ? `INH(p594) : f570;
        f570 = (f570 >= `INH(p596)) ? `INH(p596) : f570;
        f570 = (f570 > p597) ? p597 : f570;
        f571 = 4095;
        f571 = (f571 > p80) ? p80 : f571;
        f571 = (f571 >= `INH(p599)) ? `INH(p599) : f571;
        f572 = 4095;
        f572 = (f572 > p598) ? p598 : f572;
        f572 = (f572 >= `INH(p600)) ? `INH(p600) : f572;
        f573 = 4095;
        f573 = (f573 >= `INH(p80)) ? `INH(p80) : f573;
        f573 = (f573 >= `INH(p599)) ? `INH(p599) : f573;
        f573 = (f573 > p600) ? p600 : f573;
        f574 = 4095;
        f574 = (f574 >= `INH(p598)) ? `INH(p598) : f574;
        f574 = (f574 >= `INH(p600)) ? `INH(p600) : f574;
        f574 = (f574 > p601) ? p601 : f574;
        f575 = 4095;
        f575 = (f575 >= `INH(p71)) ? `INH(p71) : f575;
        f575 = (f575 > p595) ? p595 : f575;
        f575 = (f575 > p599) ? p599 : f575;
        f576 = 4095;
        f576 = (f576 > p581) ? p581 : f576;
        f576 = (f576 >= `INH(p597)) ? `INH(p597) : f576;
        f576 = (f576 >= `INH(p601)) ? `INH(p601) : f576;
        f577 = 4095;
        f577 = (f577 > p582) ? p582 : f577;
        f577 = (f577 >= `INH(p602)) ? `INH(p602) : f577;
        f578 = 4095;
        f578 = (f578 > p81) ? p81 : f578;
        f578 = (f578 >= `INH(p583)) ? `INH(p583) : f578;
        f579 = 4095;
        f579 = (f579 >= `INH(p81)) ? `INH(p81) : f579;
        f579 = (f579 >= `INH(p583)) ? `INH(p583) : f579;
        f579 = (f579 > p602) ? p602 : f579;
        f580 = 4095;
        f580 = (f580 > p72) ? p72 : f580;
        f580 = (f580 >= `INH(p582)) ? `INH(p582) : f580;
        f580 = (f580 >= `INH(p602)) ? `INH(p602) : f580;
        f581 = 4095;
        f581 = (f581 > p604) ? p604 : f581;
        f581 = (f581 >= `INH(p606)) ? `INH(p606) : f581;
        f582 = 4095;
        f582 = (f582 >= `INH(p603)) ? `INH(p603) : f582;
        f582 = (f582 >= `INH(p604)) ? `INH(p604) : f582;
        f582 = (f582 >= `INH(p606)) ? `INH(p606) : f582;
        f582 = (f582 > p607) ? p607 : f582;
        f583 = 4095;
        f583 = (f583 > p78) ? p78 : f583;
        f583 = (f583 >= `INH(p609)) ? `INH(p609) : f583;
        f584 = 4095;
        f584 = (f584 > p608) ? p608 : f584;
        f584 = (f584 >= `INH(p610)) ? `INH(p610) : f584;
        f585 = 4095;
        f585 = (f585 >= `INH(p78)) ? `INH(p78) : f585;
        f585 = (f585 >= `INH(p609)) ? `INH(p609) : f585;
        f585 = (f585 > p610) ? p610 : f585;
        f586 = 4095;
        f586 = (f586 >= `INH(p608)) ? `INH(p608) : f586;
        f586 = (f586 >= `INH(p610)) ? `INH(p610) : f586;
        f586 = (f586 > p611) ? p611 : f586;
        f587 = 4095;
        f587 = (f587 > p81) ? p81 : f587;
        f587 = (f587 >= `INH(p613)) ? `INH(p613) : f587;
        f588 = 4095;
        f588 = (f588 > p612) ? p612 : f588;
        f588 = (f588 >= `INH(p614)) ? `INH(p614) : f588;
        f589 = 4095;
        f589 = (f589 >= `INH(p81)) ? `INH(p81) : f589;
        f589 = (f589 >= `INH(p613)) ? `INH(p613) : f589;
        f589 = (f589 > p614) ? p614 : f589;
        f590 = 4095;
        f590 = (f590 >= `INH(p612)) ? `INH(p612) : f590;
        f590 = (f590 >= `INH(p614)) ? `INH(p614) : f590;
        f590 = (f590 > p615) ? p615 : f590;
        f591 = 4095;
        f591 = (f591 >= `INH(p72)) ? `INH(p72) : f591;
        f591 = (f591 > p609) ? p609 : f591;
        f591 = (f591 > p613) ? p613 : f591;
        f592 = 4095;
        f592 = (f592 > p606) ? p606 : f592;
        f592 = (f592 >= `INH(p611)) ? `INH(p611) : f592;
        f592 = (f592 >= `INH(p615)) ? `INH(p615) : f592;
        f593 = 4095;
        f593 = (f593 > p605) ? p605 : f593;
        f593 = (f593 >= `INH(p616)) ? `INH(p616) : f593;
        f594 = 4095;
        f594 = (f594 > p82) ? p82 : f594;
        f594 = (f594 >= `INH(p607)) ? `INH(p607) : f594;
        f595 = 4095;
        f595 = (f595 >= `INH(p82)) ? `INH(p82) : f595;
        f595 = (f595 >= `INH(p607)) ? `INH(p607) : f595;
        f595 = (f595 > p616) ? p616 : f595;
        f596 = 4095;
        f596 = (f596 > p73) ? p73 : f596;
        f596 = (f596 >= `INH(p605)) ? `INH(p605) : f596;
        f596 = (f596 >= `INH(p616)) ? `INH(p616) : f596;
        f597 = 4095;
        f597 = (f597 >= `INH(p618)) ? `INH(p618) : f597;
        f597 = (f597 >= `INH(p619)) ? `INH(p619) : f597;
        f597 = (f597 > p623) ? p623 : f597;
        f598 = 4095;
        f598 = (f598 > p617) ? p617 : f598;
        f598 = (f598 >= `INH(p623)) ? `INH(p623) : f598;
        f599 = 4095;
        f599 = (f599 > p621) ? p621 : f599;
        f599 = (f599 >= `INH(p623)) ? `INH(p623) : f599;
        f600 = 4095;
        f600 = (f600 >= p618/2) ? p618/2 : f600;
        f600 = (f600 >= `INH(p622)) ? `INH(p622) : f600;
        f601 = 4095;
        f601 = (f601 >= `INH(p622)) ? `INH(p622) : f601;
        f601 = (f601 > p625) ? p625 : f601;
        f602 = 4095;
        f602 = (f602 > p618) ? p618 : f602;
        f602 = (f602 >= `INH(p625)) ? `INH(p625) : f602;
        f602 = (f602 > p627) ? p627 : f602;
        f603 = 4095;
        f603 = (f603 >= `INH(p625)) ? `INH(p625) : f603;
        f603 = (f603 > p628) ? p628 : f603;
        f604 = 4095;
        f604 = (f604 > p617) ? p617 : f604;
        f604 = (f604 >= `INH(p627)) ? `INH(p627) : f604;
        f604 = (f604 >= `INH(p628)) ? `INH(p628) : f604;
        f605 = 4095;
        f605 = (f605 > p617) ? p617 : f605;
        f605 = (f605 >= `INH(p626)) ? `INH(p626) : f605;
        f605 = (f605 >= `INH(p628)) ? `INH(p628) : f605;
        f606 = 4095;
        f606 = (f606 >= `INH(p628)) ? `INH(p628) : f606;
        f606 = (f606 > p630) ? p630 : f606;
        f607 = 4095;
        f607 = (f607 > p624) ? p624 : f607;
        f607 = (f607 >= `INH(p630)) ? `INH(p630) : f607;
        f608 = 4095;
        f608 = (f608 >= `INH(p630)) ? `INH(p630) : f608;
        f608 = (f608 > p631) ? p631 : f608;
        f609 = 4095;
        f609 = (f609 > p629) ? p629 : f609;
        f609 = (f609 >= `INH(p631)) ? `INH(p631) : f609;
        f610 = 4095;
        f610 = (f610 > p619) ? p619 : f610;
        f610 = (f610 > p626) ? p626 : f610;
        f610 = (f610 >= `INH(p627)) ? `INH(p627) : f610;
        f610 = (f610 >= `INH(p631)) ? `INH(p631) : f610;
        f611 = 4095;
        f611 = (f611 > p619) ? p619 : f611;
        f611 = (f611 >= `INH(p626)) ? `INH(p626) : f611;
        f611 = (f611 >= `INH(p631)) ? `INH(p631) : f611;
        f612 = 4095;
        f612 = (f612 > p83) ? p83 : f612;
        f612 = (f612 >= `INH(p633)) ? `INH(p633) : f612;
        f613 = 4095;
        f613 = (f613 > p632) ? p632 : f613;
        f613 = (f613 >= `INH(p634)) ? `INH(p634) : f613;
        f614 = 4095;
        f614 = (f614 >= `INH(p83)) ? `INH(p83) : f614;
        f614 = (f614 >= `INH(p633)) ? `INH(p633) : f614;
        f614 = (f614 > p634) ? p634 : f614;
        f615 = 4095;
        f615 = (f615 >= `INH(p632)) ? `INH(p632) : f615;
        f615 = (f615 >= `INH(p634)) ? `INH(p634) : f615;
        f615 = (f615 > p635) ? p635 : f615;
        f616 = 4095;
        f616 = (f616 > p84) ? p84 : f616;
        f616 = (f616 >= `INH(p637)) ? `INH(p637) : f616;
        f617 = 4095;
        f617 = (f617 > p636) ? p636 : f617;
        f617 = (f617 >= `INH(p638)) ? `INH(p638) : f617;
        f618 = 4095;
        f618 = (f618 >= `INH(p84)) ? `INH(p84) : f618;
        f618 = (f618 >= `INH(p637)) ? `INH(p637) : f618;
        f618 = (f618 > p638) ? p638 : f618;
        f619 = 4095;
        f619 = (f619 >= `INH(p636)) ? `INH(p636) : f619;
        f619 = (f619 >= `INH(p638)) ? `INH(p638) : f619;
        f619 = (f619 > p639) ? p639 : f619;
        f620 = 4095;
        f620 = (f620 >= `INH(p73)) ? `INH(p73) : f620;
        f620 = (f620 > p633) ? p633 : f620;
        f620 = (f620 > p637) ? p637 : f620;
        f621 = 4095;
        f621 = (f621 > p619) ? p619 : f621;
        f621 = (f621 >= `INH(p635)) ? `INH(p635) : f621;
        f621 = (f621 >= `INH(p639)) ? `INH(p639) : f621;
        f622 = 4095;
        f622 = (f622 > p620) ? p620 : f622;
        f622 = (f622 >= `INH(p640)) ? `INH(p640) : f622;
        f623 = 4095;
        f623 = (f623 > p85) ? p85 : f623;
        f623 = (f623 >= `INH(p621)) ? `INH(p621) : f623;
        f624 = 4095;
        f624 = (f624 >= `INH(p85)) ? `INH(p85) : f624;
        f624 = (f624 >= `INH(p621)) ? `INH(p621) : f624;
        f624 = (f624 > p640) ? p640 : f624;
        f625 = 4095;
        f625 = (f625 > p74) ? p74 : f625;
        f625 = (f625 >= `INH(p620)) ? `INH(p620) : f625;
        f625 = (f625 >= `INH(p640)) ? `INH(p640) : f625;
        f626 = 4095;
        f626 = (f626 > p642) ? p642 : f626;
        f626 = (f626 >= `INH(p644)) ? `INH(p644) : f626;
        f627 = 4095;
        f627 = (f627 >= `INH(p641)) ? `INH(p641) : f627;
        f627 = (f627 >= `INH(p642)) ? `INH(p642) : f627;
        f627 = (f627 >= `INH(p644)) ? `INH(p644) : f627;
        f627 = (f627 > p645) ? p645 : f627;
        f628 = 4095;
        f628 = (f628 > p82) ? p82 : f628;
        f628 = (f628 >= `INH(p647)) ? `INH(p647) : f628;
        f629 = 4095;
        f629 = (f629 > p646) ? p646 : f629;
        f629 = (f629 >= `INH(p648)) ? `INH(p648) : f629;
        f630 = 4095;
        f630 = (f630 >= `INH(p82)) ? `INH(p82) : f630;
        f630 = (f630 >= `INH(p647)) ? `INH(p647) : f630;
        f630 = (f630 > p648) ? p648 : f630;
        f631 = 4095;
        f631 = (f631 >= `INH(p646)) ? `INH(p646) : f631;
        f631 = (f631 >= `INH(p648)) ? `INH(p648) : f631;
        f631 = (f631 > p649) ? p649 : f631;
        f632 = 4095;
        f632 = (f632 > p85) ? p85 : f632;
        f632 = (f632 >= `INH(p651)) ? `INH(p651) : f632;
        f633 = 4095;
        f633 = (f633 > p650) ? p650 : f633;
        f633 = (f633 >= `INH(p652)) ? `INH(p652) : f633;
        f634 = 4095;
        f634 = (f634 >= `INH(p85)) ? `INH(p85) : f634;
        f634 = (f634 >= `INH(p651)) ? `INH(p651) : f634;
        f634 = (f634 > p652) ? p652 : f634;
        f635 = 4095;
        f635 = (f635 >= `INH(p650)) ? `INH(p650) : f635;
        f635 = (f635 >= `INH(p652)) ? `INH(p652) : f635;
        f635 = (f635 > p653) ? p653 : f635;
        f636 = 4095;
        f636 = (f636 >= `INH(p74)) ? `INH(p74) : f636;
        f636 = (f636 > p647) ? p647 : f636;
        f636 = (f636 > p651) ? p651 : f636;
        f637 = 4095;
        f637 = (f637 > p644) ? p644 : f637;
        f637 = (f637 >= `INH(p649)) ? `INH(p649) : f637;
        f637 = (f637 >= `INH(p653)) ? `INH(p653) : f637;
        f638 = 4095;
        f638 = (f638 > p643) ? p643 : f638;
        f638 = (f638 >= `INH(p654)) ? `INH(p654) : f638;
        f639 = 4095;
        f639 = (f639 > p86) ? p86 : f639;
        f639 = (f639 >= `INH(p645)) ? `INH(p645) : f639;
        f640 = 4095;
        f640 = (f640 >= `INH(p86)) ? `INH(p86) : f640;
        f640 = (f640 >= `INH(p645)) ? `INH(p645) : f640;
        f640 = (f640 > p654) ? p654 : f640;
        f641 = 4095;
        f641 = (f641 > p75) ? p75 : f641;
        f641 = (f641 >= `INH(p643)) ? `INH(p643) : f641;
        f641 = (f641 >= `INH(p654)) ? `INH(p654) : f641;
        f642 = 4095;
        f642 = (f642 >= `INH(p656)) ? `INH(p656) : f642;
        f642 = (f642 >= `INH(p657)) ? `INH(p657) : f642;
        f642 = (f642 > p661) ? p661 : f642;
        f643 = 4095;
        f643 = (f643 > p655) ? p655 : f643;
        f643 = (f643 >= `INH(p661)) ? `INH(p661) : f643;
        f644 = 4095;
        f644 = (f644 > p659) ? p659 : f644;
        f644 = (f644 >= `INH(p661)) ? `INH(p661) : f644;
        f645 = 4095;
        f645 = (f645 >= p656/2) ? p656/2 : f645;
        f645 = (f645 >= `INH(p660)) ? `INH(p660) : f645;
        f646 = 4095;
        f646 = (f646 >= `INH(p660)) ? `INH(p660) : f646;
        f646 = (f646 > p663) ? p663 : f646;
        f647 = 4095;
        f647 = (f647 > p656) ? p656 : f647;
        f647 = (f647 >= `INH(p663)) ? `INH(p663) : f647;
        f647 = (f647 > p665) ? p665 : f647;
        f648 = 4095;
        f648 = (f648 >= `INH(p663)) ? `INH(p663) : f648;
        f648 = (f648 > p666) ? p666 : f648;
        f649 = 4095;
        f649 = (f649 > p655) ? p655 : f649;
        f649 = (f649 >= `INH(p665)) ? `INH(p665) : f649;
        f649 = (f649 >= `INH(p666)) ? `INH(p666) : f649;
        f650 = 4095;
        f650 = (f650 > p655) ? p655 : f650;
        f650 = (f650 >= `INH(p664)) ? `INH(p664) : f650;
        f650 = (f650 >= `INH(p666)) ? `INH(p666) : f650;
        f651 = 4095;
        f651 = (f651 >= `INH(p666)) ? `INH(p666) : f651;
        f651 = (f651 > p668) ? p668 : f651;
        f652 = 4095;
        f652 = (f652 > p662) ? p662 : f652;
        f652 = (f652 >= `INH(p668)) ? `INH(p668) : f652;
        f653 = 4095;
        f653 = (f653 >= `INH(p668)) ? `INH(p668) : f653;
        f653 = (f653 > p669) ? p669 : f653;
        f654 = 4095;
        f654 = (f654 > p667) ? p667 : f654;
        f654 = (f654 >= `INH(p669)) ? `INH(p669) : f654;
        f655 = 4095;
        f655 = (f655 > p657) ? p657 : f655;
        f655 = (f655 > p664) ? p664 : f655;
        f655 = (f655 >= `INH(p665)) ? `INH(p665) : f655;
        f655 = (f655 >= `INH(p669)) ? `INH(p669) : f655;
        f656 = 4095;
        f656 = (f656 > p657) ? p657 : f656;
        f656 = (f656 >= `INH(p664)) ? `INH(p664) : f656;
        f656 = (f656 >= `INH(p669)) ? `INH(p669) : f656;
        f657 = 4095;
        f657 = (f657 > p93) ? p93 : f657;
        f657 = (f657 >= `INH(p671)) ? `INH(p671) : f657;
        f658 = 4095;
        f658 = (f658 > p670) ? p670 : f658;
        f658 = (f658 >= `INH(p672)) ? `INH(p672) : f658;
        f659 = 4095;
        f659 = (f659 >= `INH(p93)) ? `INH(p93) : f659;
        f659 = (f659 >= `INH(p671)) ? `INH(p671) : f659;
        f659 = (f659 > p672) ? p672 : f659;
        f660 = 4095;
        f660 = (f660 >= `INH(p670)) ? `INH(p670) : f660;
        f660 = (f660 >= `INH(p672)) ? `INH(p672) : f660;
        f660 = (f660 > p673) ? p673 : f660;
        f661 = 4095;
        f661 = (f661 > p94) ? p94 : f661;
        f661 = (f661 >= `INH(p675)) ? `INH(p675) : f661;
        f662 = 4095;
        f662 = (f662 > p674) ? p674 : f662;
        f662 = (f662 >= `INH(p676)) ? `INH(p676) : f662;
        f663 = 4095;
        f663 = (f663 >= `INH(p94)) ? `INH(p94) : f663;
        f663 = (f663 >= `INH(p675)) ? `INH(p675) : f663;
        f663 = (f663 > p676) ? p676 : f663;
        f664 = 4095;
        f664 = (f664 >= `INH(p674)) ? `INH(p674) : f664;
        f664 = (f664 >= `INH(p676)) ? `INH(p676) : f664;
        f664 = (f664 > p677) ? p677 : f664;
        f665 = 4095;
        f665 = (f665 >= `INH(p87)) ? `INH(p87) : f665;
        f665 = (f665 > p671) ? p671 : f665;
        f665 = (f665 > p675) ? p675 : f665;
        f666 = 4095;
        f666 = (f666 > p657) ? p657 : f666;
        f666 = (f666 >= `INH(p673)) ? `INH(p673) : f666;
        f666 = (f666 >= `INH(p677)) ? `INH(p677) : f666;
        f667 = 4095;
        f667 = (f667 > p658) ? p658 : f667;
        f667 = (f667 >= `INH(p678)) ? `INH(p678) : f667;
        f668 = 4095;
        f668 = (f668 > p95) ? p95 : f668;
        f668 = (f668 >= `INH(p659)) ? `INH(p659) : f668;
        f669 = 4095;
        f669 = (f669 >= `INH(p95)) ? `INH(p95) : f669;
        f669 = (f669 >= `INH(p659)) ? `INH(p659) : f669;
        f669 = (f669 > p678) ? p678 : f669;
        f670 = 4095;
        f670 = (f670 > p88) ? p88 : f670;
        f670 = (f670 >= `INH(p658)) ? `INH(p658) : f670;
        f670 = (f670 >= `INH(p678)) ? `INH(p678) : f670;
        f671 = 4095;
        f671 = (f671 >= `INH(p680)) ? `INH(p680) : f671;
        f671 = (f671 >= `INH(p681)) ? `INH(p681) : f671;
        f671 = (f671 > p685) ? p685 : f671;
        f672 = 4095;
        f672 = (f672 > p679) ? p679 : f672;
        f672 = (f672 >= `INH(p685)) ? `INH(p685) : f672;
        f673 = 4095;
        f673 = (f673 > p683) ? p683 : f673;
        f673 = (f673 >= `INH(p685)) ? `INH(p685) : f673;
        f674 = 4095;
        f674 = (f674 >= p680/2) ? p680/2 : f674;
        f674 = (f674 >= `INH(p684)) ? `INH(p684) : f674;
        f675 = 4095;
        f675 = (f675 >= `INH(p684)) ? `INH(p684) : f675;
        f675 = (f675 > p687) ? p687 : f675;
        f676 = 4095;
        f676 = (f676 > p680) ? p680 : f676;
        f676 = (f676 >= `INH(p687)) ? `INH(p687) : f676;
        f676 = (f676 > p689) ? p689 : f676;
        f677 = 4095;
        f677 = (f677 >= `INH(p687)) ? `INH(p687) : f677;
        f677 = (f677 > p690) ? p690 : f677;
        f678 = 4095;
        f678 = (f678 > p679) ? p679 : f678;
        f678 = (f678 >= `INH(p689)) ? `INH(p689) : f678;
        f678 = (f678 >= `INH(p690)) ? `INH(p690) : f678;
        f679 = 4095;
        f679 = (f679 > p679) ? p679 : f679;
        f679 = (f679 >= `INH(p688)) ? `INH(p688) : f679;
        f679 = (f679 >= `INH(p690)) ? `INH(p690) : f679;
        f680 = 4095;
        f680 = (f680 >= `INH(p690)) ? `INH(p690) : f680;
        f680 = (f680 > p692) ? p692 : f680;
        f681 = 4095;
        f681 = (f681 > p686) ? p686 : f681;
        f681 = (f681 >= `INH(p692)) ? `INH(p692) : f681;
        f682 = 4095;
        f682 = (f682 >= `INH(p692)) ? `INH(p692) : f682;
        f682 = (f682 > p693) ? p693 : f682;
        f683 = 4095;
        f683 = (f683 > p691) ? p691 : f683;
        f683 = (f683 >= `INH(p693)) ? `INH(p693) : f683;
        f684 = 4095;
        f684 = (f684 > p681) ? p681 : f684;
        f684 = (f684 > p688) ? p688 : f684;
        f684 = (f684 >= `INH(p689)) ? `INH(p689) : f684;
        f684 = (f684 >= `INH(p693)) ? `INH(p693) : f684;
        f685 = 4095;
        f685 = (f685 > p681) ? p681 : f685;
        f685 = (f685 >= `INH(p688)) ? `INH(p688) : f685;
        f685 = (f685 >= `INH(p693)) ? `INH(p693) : f685;
        f686 = 4095;
        f686 = (f686 > p96) ? p96 : f686;
        f686 = (f686 >= `INH(p695)) ? `INH(p695) : f686;
        f687 = 4095;
        f687 = (f687 > p694) ? p694 : f687;
        f687 = (f687 >= `INH(p696)) ? `INH(p696) : f687;
        f688 = 4095;
        f688 = (f688 >= `INH(p96)) ? `INH(p96) : f688;
        f688 = (f688 >= `INH(p695)) ? `INH(p695) : f688;
        f688 = (f688 > p696) ? p696 : f688;
        f689 = 4095;
        f689 = (f689 >= `INH(p694)) ? `INH(p694) : f689;
        f689 = (f689 >= `INH(p696)) ? `INH(p696) : f689;
        f689 = (f689 > p697) ? p697 : f689;
        f690 = 4095;
        f690 = (f690 > p97) ? p97 : f690;
        f690 = (f690 >= `INH(p699)) ? `INH(p699) : f690;
        f691 = 4095;
        f691 = (f691 > p698) ? p698 : f691;
        f691 = (f691 >= `INH(p700)) ? `INH(p700) : f691;
        f692 = 4095;
        f692 = (f692 >= `INH(p97)) ? `INH(p97) : f692;
        f692 = (f692 >= `INH(p699)) ? `INH(p699) : f692;
        f692 = (f692 > p700) ? p700 : f692;
        f693 = 4095;
        f693 = (f693 >= `INH(p698)) ? `INH(p698) : f693;
        f693 = (f693 >= `INH(p700)) ? `INH(p700) : f693;
        f693 = (f693 > p701) ? p701 : f693;
        f694 = 4095;
        f694 = (f694 >= `INH(p88)) ? `INH(p88) : f694;
        f694 = (f694 > p695) ? p695 : f694;
        f694 = (f694 > p699) ? p699 : f694;
        f695 = 4095;
        f695 = (f695 > p681) ? p681 : f695;
        f695 = (f695 >= `INH(p697)) ? `INH(p697) : f695;
        f695 = (f695 >= `INH(p701)) ? `INH(p701) : f695;
        f696 = 4095;
        f696 = (f696 > p682) ? p682 : f696;
        f696 = (f696 >= `INH(p702)) ? `INH(p702) : f696;
        f697 = 4095;
        f697 = (f697 > p98) ? p98 : f697;
        f697 = (f697 >= `INH(p683)) ? `INH(p683) : f697;
        f698 = 4095;
        f698 = (f698 >= `INH(p98)) ? `INH(p98) : f698;
        f698 = (f698 >= `INH(p683)) ? `INH(p683) : f698;
        f698 = (f698 > p702) ? p702 : f698;
        f699 = 4095;
        f699 = (f699 > p89) ? p89 : f699;
        f699 = (f699 >= `INH(p682)) ? `INH(p682) : f699;
        f699 = (f699 >= `INH(p702)) ? `INH(p702) : f699;
        f700 = 4095;
        f700 = (f700 > p704) ? p704 : f700;
        f700 = (f700 >= `INH(p706)) ? `INH(p706) : f700;
        f701 = 4095;
        f701 = (f701 >= `INH(p703)) ? `INH(p703) : f701;
        f701 = (f701 >= `INH(p704)) ? `INH(p704) : f701;
        f701 = (f701 >= `INH(p706)) ? `INH(p706) : f701;
        f701 = (f701 > p707) ? p707 : f701;
        f702 = 4095;
        f702 = (f702 > p95) ? p95 : f702;
        f702 = (f702 >= `INH(p709)) ? `INH(p709) : f702;
        f703 = 4095;
        f703 = (f703 > p708) ? p708 : f703;
        f703 = (f703 >= `INH(p710)) ? `INH(p710) : f703;
        f704 = 4095;
        f704 = (f704 >= `INH(p95)) ? `INH(p95) : f704;
        f704 = (f704 >= `INH(p709)) ? `INH(p709) : f704;
        f704 = (f704 > p710) ? p710 : f704;
        f705 = 4095;
        f705 = (f705 >= `INH(p708)) ? `INH(p708) : f705;
        f705 = (f705 >= `INH(p710)) ? `INH(p710) : f705;
        f705 = (f705 > p711) ? p711 : f705;
        f706 = 4095;
        f706 = (f706 > p98) ? p98 : f706;
        f706 = (f706 >= `INH(p713)) ? `INH(p713) : f706;
        f707 = 4095;
        f707 = (f707 > p712) ? p712 : f707;
        f707 = (f707 >= `INH(p714)) ? `INH(p714) : f707;
        f708 = 4095;
        f708 = (f708 >= `INH(p98)) ? `INH(p98) : f708;
        f708 = (f708 >= `INH(p713)) ? `INH(p713) : f708;
        f708 = (f708 > p714) ? p714 : f708;
        f709 = 4095;
        f709 = (f709 >= `INH(p712)) ? `INH(p712) : f709;
        f709 = (f709 >= `INH(p714)) ? `INH(p714) : f709;
        f709 = (f709 > p715) ? p715 : f709;
        f710 = 4095;
        f710 = (f710 >= `INH(p89)) ? `INH(p89) : f710;
        f710 = (f710 > p709) ? p709 : f710;
        f710 = (f710 > p713) ? p713 : f710;
        f711 = 4095;
        f711 = (f711 > p706) ? p706 : f711;
        f711 = (f711 >= `INH(p711)) ? `INH(p711) : f711;
        f711 = (f711 >= `INH(p715)) ? `INH(p715) : f711;
        f712 = 4095;
        f712 = (f712 > p705) ? p705 : f712;
        f712 = (f712 >= `INH(p716)) ? `INH(p716) : f712;
        f713 = 4095;
        f713 = (f713 > p99) ? p99 : f713;
        f713 = (f713 >= `INH(p707)) ? `INH(p707) : f713;
        f714 = 4095;
        f714 = (f714 >= `INH(p99)) ? `INH(p99) : f714;
        f714 = (f714 >= `INH(p707)) ? `INH(p707) : f714;
        f714 = (f714 > p716) ? p716 : f714;
        f715 = 4095;
        f715 = (f715 > p90) ? p90 : f715;
        f715 = (f715 >= `INH(p705)) ? `INH(p705) : f715;
        f715 = (f715 >= `INH(p716)) ? `INH(p716) : f715;
        f716 = 4095;
        f716 = (f716 >= `INH(p718)) ? `INH(p718) : f716;
        f716 = (f716 >= `INH(p719)) ? `INH(p719) : f716;
        f716 = (f716 > p723) ? p723 : f716;
        f717 = 4095;
        f717 = (f717 > p717) ? p717 : f717;
        f717 = (f717 >= `INH(p723)) ? `INH(p723) : f717;
        f718 = 4095;
        f718 = (f718 > p721) ? p721 : f718;
        f718 = (f718 >= `INH(p723)) ? `INH(p723) : f718;
        f719 = 4095;
        f719 = (f719 >= p718/2) ? p718/2 : f719;
        f719 = (f719 >= `INH(p722)) ? `INH(p722) : f719;
        f720 = 4095;
        f720 = (f720 >= `INH(p722)) ? `INH(p722) : f720;
        f720 = (f720 > p725) ? p725 : f720;
        f721 = 4095;
        f721 = (f721 > p718) ? p718 : f721;
        f721 = (f721 >= `INH(p725)) ? `INH(p725) : f721;
        f721 = (f721 > p727) ? p727 : f721;
        f722 = 4095;
        f722 = (f722 >= `INH(p725)) ? `INH(p725) : f722;
        f722 = (f722 > p728) ? p728 : f722;
        f723 = 4095;
        f723 = (f723 > p717) ? p717 : f723;
        f723 = (f723 >= `INH(p727)) ? `INH(p727) : f723;
        f723 = (f723 >= `INH(p728)) ? `INH(p728) : f723;
        f724 = 4095;
        f724 = (f724 > p717) ? p717 : f724;
        f724 = (f724 >= `INH(p726)) ? `INH(p726) : f724;
        f724 = (f724 >= `INH(p728)) ? `INH(p728) : f724;
        f725 = 4095;
        f725 = (f725 >= `INH(p728)) ? `INH(p728) : f725;
        f725 = (f725 > p730) ? p730 : f725;
        f726 = 4095;
        f726 = (f726 > p724) ? p724 : f726;
        f726 = (f726 >= `INH(p730)) ? `INH(p730) : f726;
        f727 = 4095;
        f727 = (f727 >= `INH(p730)) ? `INH(p730) : f727;
        f727 = (f727 > p731) ? p731 : f727;
        f728 = 4095;
        f728 = (f728 > p729) ? p729 : f728;
        f728 = (f728 >= `INH(p731)) ? `INH(p731) : f728;
        f729 = 4095;
        f729 = (f729 > p719) ? p719 : f729;
        f729 = (f729 > p726) ? p726 : f729;
        f729 = (f729 >= `INH(p727)) ? `INH(p727) : f729;
        f729 = (f729 >= `INH(p731)) ? `INH(p731) : f729;
        f730 = 4095;
        f730 = (f730 > p719) ? p719 : f730;
        f730 = (f730 >= `INH(p726)) ? `INH(p726) : f730;
        f730 = (f730 >= `INH(p731)) ? `INH(p731) : f730;
        f731 = 4095;
        f731 = (f731 > p100) ? p100 : f731;
        f731 = (f731 >= `INH(p733)) ? `INH(p733) : f731;
        f732 = 4095;
        f732 = (f732 > p732) ? p732 : f732;
        f732 = (f732 >= `INH(p734)) ? `INH(p734) : f732;
        f733 = 4095;
        f733 = (f733 >= `INH(p100)) ? `INH(p100) : f733;
        f733 = (f733 >= `INH(p733)) ? `INH(p733) : f733;
        f733 = (f733 > p734) ? p734 : f733;
        f734 = 4095;
        f734 = (f734 >= `INH(p732)) ? `INH(p732) : f734;
        f734 = (f734 >= `INH(p734)) ? `INH(p734) : f734;
        f734 = (f734 > p735) ? p735 : f734;
        f735 = 4095;
        f735 = (f735 > p101) ? p101 : f735;
        f735 = (f735 >= `INH(p737)) ? `INH(p737) : f735;
        f736 = 4095;
        f736 = (f736 > p736) ? p736 : f736;
        f736 = (f736 >= `INH(p738)) ? `INH(p738) : f736;
        f737 = 4095;
        f737 = (f737 >= `INH(p101)) ? `INH(p101) : f737;
        f737 = (f737 >= `INH(p737)) ? `INH(p737) : f737;
        f737 = (f737 > p738) ? p738 : f737;
        f738 = 4095;
        f738 = (f738 >= `INH(p736)) ? `INH(p736) : f738;
        f738 = (f738 >= `INH(p738)) ? `INH(p738) : f738;
        f738 = (f738 > p739) ? p739 : f738;
        f739 = 4095;
        f739 = (f739 >= `INH(p90)) ? `INH(p90) : f739;
        f739 = (f739 > p733) ? p733 : f739;
        f739 = (f739 > p737) ? p737 : f739;
        f740 = 4095;
        f740 = (f740 > p719) ? p719 : f740;
        f740 = (f740 >= `INH(p735)) ? `INH(p735) : f740;
        f740 = (f740 >= `INH(p739)) ? `INH(p739) : f740;
        f741 = 4095;
        f741 = (f741 > p720) ? p720 : f741;
        f741 = (f741 >= `INH(p740)) ? `INH(p740) : f741;
        f742 = 4095;
        f742 = (f742 > p102) ? p102 : f742;
        f742 = (f742 >= `INH(p721)) ? `INH(p721) : f742;
        f743 = 4095;
        f743 = (f743 >= `INH(p102)) ? `INH(p102) : f743;
        f743 = (f743 >= `INH(p721)) ? `INH(p721) : f743;
        f743 = (f743 > p740) ? p740 : f743;
        f744 = 4095;
        f744 = (f744 > p91) ? p91 : f744;
        f744 = (f744 >= `INH(p720)) ? `INH(p720) : f744;
        f744 = (f744 >= `INH(p740)) ? `INH(p740) : f744;
        f745 = 4095;
        f745 = (f745 > p742) ? p742 : f745;
        f745 = (f745 >= `INH(p744)) ? `INH(p744) : f745;
        f746 = 4095;
        f746 = (f746 >= `INH(p741)) ? `INH(p741) : f746;
        f746 = (f746 >= `INH(p742)) ? `INH(p742) : f746;
        f746 = (f746 >= `INH(p744)) ? `INH(p744) : f746;
        f746 = (f746 > p745) ? p745 : f746;
        f747 = 4095;
        f747 = (f747 > p99) ? p99 : f747;
        f747 = (f747 >= `INH(p747)) ? `INH(p747) : f747;
        f748 = 4095;
        f748 = (f748 > p746) ? p746 : f748;
        f748 = (f748 >= `INH(p748)) ? `INH(p748) : f748;
        f749 = 4095;
        f749 = (f749 >= `INH(p99)) ? `INH(p99) : f749;
        f749 = (f749 >= `INH(p747)) ? `INH(p747) : f749;
        f749 = (f749 > p748) ? p748 : f749;
        f750 = 4095;
        f750 = (f750 >= `INH(p746)) ? `INH(p746) : f750;
        f750 = (f750 >= `INH(p748)) ? `INH(p748) : f750;
        f750 = (f750 > p749) ? p749 : f750;
        f751 = 4095;
        f751 = (f751 > p102) ? p102 : f751;
        f751 = (f751 >= `INH(p751)) ? `INH(p751) : f751;
        f752 = 4095;
        f752 = (f752 > p750) ? p750 : f752;
        f752 = (f752 >= `INH(p752)) ? `INH(p752) : f752;
        f753 = 4095;
        f753 = (f753 >= `INH(p102)) ? `INH(p102) : f753;
        f753 = (f753 >= `INH(p751)) ? `INH(p751) : f753;
        f753 = (f753 > p752) ? p752 : f753;
        f754 = 4095;
        f754 = (f754 >= `INH(p750)) ? `INH(p750) : f754;
        f754 = (f754 >= `INH(p752)) ? `INH(p752) : f754;
        f754 = (f754 > p753) ? p753 : f754;
        f755 = 4095;
        f755 = (f755 >= `INH(p91)) ? `INH(p91) : f755;
        f755 = (f755 > p747) ? p747 : f755;
        f755 = (f755 > p751) ? p751 : f755;
        f756 = 4095;
        f756 = (f756 > p744) ? p744 : f756;
        f756 = (f756 >= `INH(p749)) ? `INH(p749) : f756;
        f756 = (f756 >= `INH(p753)) ? `INH(p753) : f756;
        f757 = 4095;
        f757 = (f757 > p743) ? p743 : f757;
        f757 = (f757 >= `INH(p754)) ? `INH(p754) : f757;
        f758 = 4095;
        f758 = (f758 > p103) ? p103 : f758;
        f758 = (f758 >= `INH(p745)) ? `INH(p745) : f758;
        f759 = 4095;
        f759 = (f759 >= `INH(p103)) ? `INH(p103) : f759;
        f759 = (f759 >= `INH(p745)) ? `INH(p745) : f759;
        f759 = (f759 > p754) ? p754 : f759;
        f760 = 4095;
        f760 = (f760 > p92) ? p92 : f760;
        f760 = (f760 >= `INH(p743)) ? `INH(p743) : f760;
        f760 = (f760 >= `INH(p754)) ? `INH(p754) : f760;
        f761 = 4095;
        f761 = (f761 >= `INH(p756)) ? `INH(p756) : f761;
        f761 = (f761 >= `INH(p757)) ? `INH(p757) : f761;
        f761 = (f761 > p761) ? p761 : f761;
        f762 = 4095;
        f762 = (f762 > p755) ? p755 : f762;
        f762 = (f762 >= `INH(p761)) ? `INH(p761) : f762;
        f763 = 4095;
        f763 = (f763 > p759) ? p759 : f763;
        f763 = (f763 >= `INH(p761)) ? `INH(p761) : f763;
        f764 = 4095;
        f764 = (f764 >= p756/2) ? p756/2 : f764;
        f764 = (f764 >= `INH(p760)) ? `INH(p760) : f764;
        f765 = 4095;
        f765 = (f765 >= `INH(p760)) ? `INH(p760) : f765;
        f765 = (f765 > p763) ? p763 : f765;
        f766 = 4095;
        f766 = (f766 > p756) ? p756 : f766;
        f766 = (f766 >= `INH(p763)) ? `INH(p763) : f766;
        f766 = (f766 > p765) ? p765 : f766;
        f767 = 4095;
        f767 = (f767 >= `INH(p763)) ? `INH(p763) : f767;
        f767 = (f767 > p766) ? p766 : f767;
        f768 = 4095;
        f768 = (f768 > p755) ? p755 : f768;
        f768 = (f768 >= `INH(p765)) ? `INH(p765) : f768;
        f768 = (f768 >= `INH(p766)) ? `INH(p766) : f768;
        f769 = 4095;
        f769 = (f769 > p755) ? p755 : f769;
        f769 = (f769 >= `INH(p764)) ? `INH(p764) : f769;
        f769 = (f769 >= `INH(p766)) ? `INH(p766) : f769;
        f770 = 4095;
        f770 = (f770 >= `INH(p766)) ? `INH(p766) : f770;
        f770 = (f770 > p768) ? p768 : f770;
        f771 = 4095;
        f771 = (f771 > p762) ? p762 : f771;
        f771 = (f771 >= `INH(p768)) ? `INH(p768) : f771;
        f772 = 4095;
        f772 = (f772 >= `INH(p768)) ? `INH(p768) : f772;
        f772 = (f772 > p769) ? p769 : f772;
        f773 = 4095;
        f773 = (f773 > p767) ? p767 : f773;
        f773 = (f773 >= `INH(p769)) ? `INH(p769) : f773;
        f774 = 4095;
        f774 = (f774 > p757) ? p757 : f774;
        f774 = (f774 > p764) ? p764 : f774;
        f774 = (f774 >= `INH(p765)) ? `INH(p765) : f774;
        f774 = (f774 >= `INH(p769)) ? `INH(p769) : f774;
        f775 = 4095;
        f775 = (f775 > p757) ? p757 : f775;
        f775 = (f775 >= `INH(p764)) ? `INH(p764) : f775;
        f775 = (f775 >= `INH(p769)) ? `INH(p769) : f775;
        f776 = 4095;
        f776 = (f776 > p110) ? p110 : f776;
        f776 = (f776 >= `INH(p771)) ? `INH(p771) : f776;
        f777 = 4095;
        f777 = (f777 > p770) ? p770 : f777;
        f777 = (f777 >= `INH(p772)) ? `INH(p772) : f777;
        f778 = 4095;
        f778 = (f778 >= `INH(p110)) ? `INH(p110) : f778;
        f778 = (f778 >= `INH(p771)) ? `INH(p771) : f778;
        f778 = (f778 > p772) ? p772 : f778;
        f779 = 4095;
        f779 = (f779 >= `INH(p770)) ? `INH(p770) : f779;
        f779 = (f779 >= `INH(p772)) ? `INH(p772) : f779;
        f779 = (f779 > p773) ? p773 : f779;
        f780 = 4095;
        f780 = (f780 > p111) ? p111 : f780;
        f780 = (f780 >= `INH(p775)) ? `INH(p775) : f780;
        f781 = 4095;
        f781 = (f781 > p774) ? p774 : f781;
        f781 = (f781 >= `INH(p776)) ? `INH(p776) : f781;
        f782 = 4095;
        f782 = (f782 >= `INH(p111)) ? `INH(p111) : f782;
        f782 = (f782 >= `INH(p775)) ? `INH(p775) : f782;
        f782 = (f782 > p776) ? p776 : f782;
        f783 = 4095;
        f783 = (f783 >= `INH(p774)) ? `INH(p774) : f783;
        f783 = (f783 >= `INH(p776)) ? `INH(p776) : f783;
        f783 = (f783 > p777) ? p777 : f783;
        f784 = 4095;
        f784 = (f784 >= `INH(p104)) ? `INH(p104) : f784;
        f784 = (f784 > p771) ? p771 : f784;
        f784 = (f784 > p775) ? p775 : f784;
        f785 = 4095;
        f785 = (f785 > p757) ? p757 : f785;
        f785 = (f785 >= `INH(p773)) ? `INH(p773) : f785;
        f785 = (f785 >= `INH(p777)) ? `INH(p777) : f785;
        f786 = 4095;
        f786 = (f786 > p758) ? p758 : f786;
        f786 = (f786 >= `INH(p778)) ? `INH(p778) : f786;
        f787 = 4095;
        f787 = (f787 > p112) ? p112 : f787;
        f787 = (f787 >= `INH(p759)) ? `INH(p759) : f787;
        f788 = 4095;
        f788 = (f788 >= `INH(p112)) ? `INH(p112) : f788;
        f788 = (f788 >= `INH(p759)) ? `INH(p759) : f788;
        f788 = (f788 > p778) ? p778 : f788;
        f789 = 4095;
        f789 = (f789 > p105) ? p105 : f789;
        f789 = (f789 >= `INH(p758)) ? `INH(p758) : f789;
        f789 = (f789 >= `INH(p778)) ? `INH(p778) : f789;
        f790 = 4095;
        f790 = (f790 >= `INH(p780)) ? `INH(p780) : f790;
        f790 = (f790 >= `INH(p781)) ? `INH(p781) : f790;
        f790 = (f790 > p785) ? p785 : f790;
        f791 = 4095;
        f791 = (f791 > p779) ? p779 : f791;
        f791 = (f791 >= `INH(p785)) ? `INH(p785) : f791;
        f792 = 4095;
        f792 = (f792 > p783) ? p783 : f792;
        f792 = (f792 >= `INH(p785)) ? `INH(p785) : f792;
        f793 = 4095;
        f793 = (f793 >= p780/2) ? p780/2 : f793;
        f793 = (f793 >= `INH(p784)) ? `INH(p784) : f793;
        f794 = 4095;
        f794 = (f794 >= `INH(p784)) ? `INH(p784) : f794;
        f794 = (f794 > p787) ? p787 : f794;
        f795 = 4095;
        f795 = (f795 > p780) ? p780 : f795;
        f795 = (f795 >= `INH(p787)) ? `INH(p787) : f795;
        f795 = (f795 > p789) ? p789 : f795;
        f796 = 4095;
        f796 = (f796 >= `INH(p787)) ? `INH(p787) : f796;
        f796 = (f796 > p790) ? p790 : f796;
        f797 = 4095;
        f797 = (f797 > p779) ? p779 : f797;
        f797 = (f797 >= `INH(p789)) ? `INH(p789) : f797;
        f797 = (f797 >= `INH(p790)) ? `INH(p790) : f797;
        f798 = 4095;
        f798 = (f798 > p779) ? p779 : f798;
        f798 = (f798 >= `INH(p788)) ? `INH(p788) : f798;
        f798 = (f798 >= `INH(p790)) ? `INH(p790) : f798;
        f799 = 4095;
        f799 = (f799 >= `INH(p790)) ? `INH(p790) : f799;
        f799 = (f799 > p792) ? p792 : f799;
        f800 = 4095;
        f800 = (f800 > p786) ? p786 : f800;
        f800 = (f800 >= `INH(p792)) ? `INH(p792) : f800;
        f801 = 4095;
        f801 = (f801 >= `INH(p792)) ? `INH(p792) : f801;
        f801 = (f801 > p793) ? p793 : f801;
        f802 = 4095;
        f802 = (f802 > p791) ? p791 : f802;
        f802 = (f802 >= `INH(p793)) ? `INH(p793) : f802;
        f803 = 4095;
        f803 = (f803 > p781) ? p781 : f803;
        f803 = (f803 > p788) ? p788 : f803;
        f803 = (f803 >= `INH(p789)) ? `INH(p789) : f803;
        f803 = (f803 >= `INH(p793)) ? `INH(p793) : f803;
        f804 = 4095;
        f804 = (f804 > p781) ? p781 : f804;
        f804 = (f804 >= `INH(p788)) ? `INH(p788) : f804;
        f804 = (f804 >= `INH(p793)) ? `INH(p793) : f804;
        f805 = 4095;
        f805 = (f805 > p113) ? p113 : f805;
        f805 = (f805 >= `INH(p795)) ? `INH(p795) : f805;
        f806 = 4095;
        f806 = (f806 > p794) ? p794 : f806;
        f806 = (f806 >= `INH(p796)) ? `INH(p796) : f806;
        f807 = 4095;
        f807 = (f807 >= `INH(p113)) ? `INH(p113) : f807;
        f807 = (f807 >= `INH(p795)) ? `INH(p795) : f807;
        f807 = (f807 > p796) ? p796 : f807;
        f808 = 4095;
        f808 = (f808 >= `INH(p794)) ? `INH(p794) : f808;
        f808 = (f808 >= `INH(p796)) ? `INH(p796) : f808;
        f808 = (f808 > p797) ? p797 : f808;
        f809 = 4095;
        f809 = (f809 > p114) ? p114 : f809;
        f809 = (f809 >= `INH(p799)) ? `INH(p799) : f809;
        f810 = 4095;
        f810 = (f810 > p798) ? p798 : f810;
        f810 = (f810 >= `INH(p800)) ? `INH(p800) : f810;
        f811 = 4095;
        f811 = (f811 >= `INH(p114)) ? `INH(p114) : f811;
        f811 = (f811 >= `INH(p799)) ? `INH(p799) : f811;
        f811 = (f811 > p800) ? p800 : f811;
        f812 = 4095;
        f812 = (f812 >= `INH(p798)) ? `INH(p798) : f812;
        f812 = (f812 >= `INH(p800)) ? `INH(p800) : f812;
        f812 = (f812 > p801) ? p801 : f812;
        f813 = 4095;
        f813 = (f813 >= `INH(p105)) ? `INH(p105) : f813;
        f813 = (f813 > p795) ? p795 : f813;
        f813 = (f813 > p799) ? p799 : f813;
        f814 = 4095;
        f814 = (f814 > p781) ? p781 : f814;
        f814 = (f814 >= `INH(p797)) ? `INH(p797) : f814;
        f814 = (f814 >= `INH(p801)) ? `INH(p801) : f814;
        f815 = 4095;
        f815 = (f815 > p782) ? p782 : f815;
        f815 = (f815 >= `INH(p802)) ? `INH(p802) : f815;
        f816 = 4095;
        f816 = (f816 > p115) ? p115 : f816;
        f816 = (f816 >= `INH(p783)) ? `INH(p783) : f816;
        f817 = 4095;
        f817 = (f817 >= `INH(p115)) ? `INH(p115) : f817;
        f817 = (f817 >= `INH(p783)) ? `INH(p783) : f817;
        f817 = (f817 > p802) ? p802 : f817;
        f818 = 4095;
        f818 = (f818 > p106) ? p106 : f818;
        f818 = (f818 >= `INH(p782)) ? `INH(p782) : f818;
        f818 = (f818 >= `INH(p802)) ? `INH(p802) : f818;
        f819 = 4095;
        f819 = (f819 > p804) ? p804 : f819;
        f819 = (f819 >= `INH(p806)) ? `INH(p806) : f819;
        f820 = 4095;
        f820 = (f820 >= `INH(p803)) ? `INH(p803) : f820;
        f820 = (f820 >= `INH(p804)) ? `INH(p804) : f820;
        f820 = (f820 >= `INH(p806)) ? `INH(p806) : f820;
        f820 = (f820 > p807) ? p807 : f820;
        f821 = 4095;
        f821 = (f821 > p112) ? p112 : f821;
        f821 = (f821 >= `INH(p809)) ? `INH(p809) : f821;
        f822 = 4095;
        f822 = (f822 > p808) ? p808 : f822;
        f822 = (f822 >= `INH(p810)) ? `INH(p810) : f822;
        f823 = 4095;
        f823 = (f823 >= `INH(p112)) ? `INH(p112) : f823;
        f823 = (f823 >= `INH(p809)) ? `INH(p809) : f823;
        f823 = (f823 > p810) ? p810 : f823;
        f824 = 4095;
        f824 = (f824 >= `INH(p808)) ? `INH(p808) : f824;
        f824 = (f824 >= `INH(p810)) ? `INH(p810) : f824;
        f824 = (f824 > p811) ? p811 : f824;
        f825 = 4095;
        f825 = (f825 > p115) ? p115 : f825;
        f825 = (f825 >= `INH(p813)) ? `INH(p813) : f825;
        f826 = 4095;
        f826 = (f826 > p812) ? p812 : f826;
        f826 = (f826 >= `INH(p814)) ? `INH(p814) : f826;
        f827 = 4095;
        f827 = (f827 >= `INH(p115)) ? `INH(p115) : f827;
        f827 = (f827 >= `INH(p813)) ? `INH(p813) : f827;
        f827 = (f827 > p814) ? p814 : f827;
        f828 = 4095;
        f828 = (f828 >= `INH(p812)) ? `INH(p812) : f828;
        f828 = (f828 >= `INH(p814)) ? `INH(p814) : f828;
        f828 = (f828 > p815) ? p815 : f828;
        f829 = 4095;
        f829 = (f829 >= `INH(p106)) ? `INH(p106) : f829;
        f829 = (f829 > p809) ? p809 : f829;
        f829 = (f829 > p813) ? p813 : f829;
        f830 = 4095;
        f830 = (f830 > p806) ? p806 : f830;
        f830 = (f830 >= `INH(p811)) ? `INH(p811) : f830;
        f830 = (f830 >= `INH(p815)) ? `INH(p815) : f830;
        f831 = 4095;
        f831 = (f831 > p805) ? p805 : f831;
        f831 = (f831 >= `INH(p816)) ? `INH(p816) : f831;
        f832 = 4095;
        f832 = (f832 > p116) ? p116 : f832;
        f832 = (f832 >= `INH(p807)) ? `INH(p807) : f832;
        f833 = 4095;
        f833 = (f833 >= `INH(p116)) ? `INH(p116) : f833;
        f833 = (f833 >= `INH(p807)) ? `INH(p807) : f833;
        f833 = (f833 > p816) ? p816 : f833;
        f834 = 4095;
        f834 = (f834 > p107) ? p107 : f834;
        f834 = (f834 >= `INH(p805)) ? `INH(p805) : f834;
        f834 = (f834 >= `INH(p816)) ? `INH(p816) : f834;
        f835 = 4095;
        f835 = (f835 >= `INH(p818)) ? `INH(p818) : f835;
        f835 = (f835 >= `INH(p819)) ? `INH(p819) : f835;
        f835 = (f835 > p823) ? p823 : f835;
        f836 = 4095;
        f836 = (f836 > p817) ? p817 : f836;
        f836 = (f836 >= `INH(p823)) ? `INH(p823) : f836;
        f837 = 4095;
        f837 = (f837 > p821) ? p821 : f837;
        f837 = (f837 >= `INH(p823)) ? `INH(p823) : f837;
        f838 = 4095;
        f838 = (f838 >= p818/2) ? p818/2 : f838;
        f838 = (f838 >= `INH(p822)) ? `INH(p822) : f838;
        f839 = 4095;
        f839 = (f839 >= `INH(p822)) ? `INH(p822) : f839;
        f839 = (f839 > p825) ? p825 : f839;
        f840 = 4095;
        f840 = (f840 > p818) ? p818 : f840;
        f840 = (f840 >= `INH(p825)) ? `INH(p825) : f840;
        f840 = (f840 > p827) ? p827 : f840;
        f841 = 4095;
        f841 = (f841 >= `INH(p825)) ? `INH(p825) : f841;
        f841 = (f841 > p828) ? p828 : f841;
        f842 = 4095;
        f842 = (f842 > p817) ? p817 : f842;
        f842 = (f842 >= `INH(p827)) ? `INH(p827) : f842;
        f842 = (f842 >= `INH(p828)) ? `INH(p828) : f842;
        f843 = 4095;
        f843 = (f843 > p817) ? p817 : f843;
        f843 = (f843 >= `INH(p826)) ? `INH(p826) : f843;
        f843 = (f843 >= `INH(p828)) ? `INH(p828) : f843;
        f844 = 4095;
        f844 = (f844 >= `INH(p828)) ? `INH(p828) : f844;
        f844 = (f844 > p830) ? p830 : f844;
        f845 = 4095;
        f845 = (f845 > p824) ? p824 : f845;
        f845 = (f845 >= `INH(p830)) ? `INH(p830) : f845;
        f846 = 4095;
        f846 = (f846 >= `INH(p830)) ? `INH(p830) : f846;
        f846 = (f846 > p831) ? p831 : f846;
        f847 = 4095;
        f847 = (f847 > p829) ? p829 : f847;
        f847 = (f847 >= `INH(p831)) ? `INH(p831) : f847;
        f848 = 4095;
        f848 = (f848 > p819) ? p819 : f848;
        f848 = (f848 > p826) ? p826 : f848;
        f848 = (f848 >= `INH(p827)) ? `INH(p827) : f848;
        f848 = (f848 >= `INH(p831)) ? `INH(p831) : f848;
        f849 = 4095;
        f849 = (f849 > p819) ? p819 : f849;
        f849 = (f849 >= `INH(p826)) ? `INH(p826) : f849;
        f849 = (f849 >= `INH(p831)) ? `INH(p831) : f849;
        f850 = 4095;
        f850 = (f850 > p117) ? p117 : f850;
        f850 = (f850 >= `INH(p833)) ? `INH(p833) : f850;
        f851 = 4095;
        f851 = (f851 > p832) ? p832 : f851;
        f851 = (f851 >= `INH(p834)) ? `INH(p834) : f851;
        f852 = 4095;
        f852 = (f852 >= `INH(p117)) ? `INH(p117) : f852;
        f852 = (f852 >= `INH(p833)) ? `INH(p833) : f852;
        f852 = (f852 > p834) ? p834 : f852;
        f853 = 4095;
        f853 = (f853 >= `INH(p832)) ? `INH(p832) : f853;
        f853 = (f853 >= `INH(p834)) ? `INH(p834) : f853;
        f853 = (f853 > p835) ? p835 : f853;
        f854 = 4095;
        f854 = (f854 > p118) ? p118 : f854;
        f854 = (f854 >= `INH(p837)) ? `INH(p837) : f854;
        f855 = 4095;
        f855 = (f855 > p836) ? p836 : f855;
        f855 = (f855 >= `INH(p838)) ? `INH(p838) : f855;
        f856 = 4095;
        f856 = (f856 >= `INH(p118)) ? `INH(p118) : f856;
        f856 = (f856 >= `INH(p837)) ? `INH(p837) : f856;
        f856 = (f856 > p838) ? p838 : f856;
        f857 = 4095;
        f857 = (f857 >= `INH(p836)) ? `INH(p836) : f857;
        f857 = (f857 >= `INH(p838)) ? `INH(p838) : f857;
        f857 = (f857 > p839) ? p839 : f857;
        f858 = 4095;
        f858 = (f858 >= `INH(p107)) ? `INH(p107) : f858;
        f858 = (f858 > p833) ? p833 : f858;
        f858 = (f858 > p837) ? p837 : f858;
        f859 = 4095;
        f859 = (f859 > p819) ? p819 : f859;
        f859 = (f859 >= `INH(p835)) ? `INH(p835) : f859;
        f859 = (f859 >= `INH(p839)) ? `INH(p839) : f859;
        f860 = 4095;
        f860 = (f860 > p820) ? p820 : f860;
        f860 = (f860 >= `INH(p840)) ? `INH(p840) : f860;
        f861 = 4095;
        f861 = (f861 > p119) ? p119 : f861;
        f861 = (f861 >= `INH(p821)) ? `INH(p821) : f861;
        f862 = 4095;
        f862 = (f862 >= `INH(p119)) ? `INH(p119) : f862;
        f862 = (f862 >= `INH(p821)) ? `INH(p821) : f862;
        f862 = (f862 > p840) ? p840 : f862;
        f863 = 4095;
        f863 = (f863 > p108) ? p108 : f863;
        f863 = (f863 >= `INH(p820)) ? `INH(p820) : f863;
        f863 = (f863 >= `INH(p840)) ? `INH(p840) : f863;
        f864 = 4095;
        f864 = (f864 > p842) ? p842 : f864;
        f864 = (f864 >= `INH(p844)) ? `INH(p844) : f864;
        f865 = 4095;
        f865 = (f865 >= `INH(p841)) ? `INH(p841) : f865;
        f865 = (f865 >= `INH(p842)) ? `INH(p842) : f865;
        f865 = (f865 >= `INH(p844)) ? `INH(p844) : f865;
        f865 = (f865 > p845) ? p845 : f865;
        f866 = 4095;
        f866 = (f866 > p116) ? p116 : f866;
        f866 = (f866 >= `INH(p847)) ? `INH(p847) : f866;
        f867 = 4095;
        f867 = (f867 > p846) ? p846 : f867;
        f867 = (f867 >= `INH(p848)) ? `INH(p848) : f867;
        f868 = 4095;
        f868 = (f868 >= `INH(p116)) ? `INH(p116) : f868;
        f868 = (f868 >= `INH(p847)) ? `INH(p847) : f868;
        f868 = (f868 > p848) ? p848 : f868;
        f869 = 4095;
        f869 = (f869 >= `INH(p846)) ? `INH(p846) : f869;
        f869 = (f869 >= `INH(p848)) ? `INH(p848) : f869;
        f869 = (f869 > p849) ? p849 : f869;
        f870 = 4095;
        f870 = (f870 > p119) ? p119 : f870;
        f870 = (f870 >= `INH(p851)) ? `INH(p851) : f870;
        f871 = 4095;
        f871 = (f871 > p850) ? p850 : f871;
        f871 = (f871 >= `INH(p852)) ? `INH(p852) : f871;
        f872 = 4095;
        f872 = (f872 >= `INH(p119)) ? `INH(p119) : f872;
        f872 = (f872 >= `INH(p851)) ? `INH(p851) : f872;
        f872 = (f872 > p852) ? p852 : f872;
        f873 = 4095;
        f873 = (f873 >= `INH(p850)) ? `INH(p850) : f873;
        f873 = (f873 >= `INH(p852)) ? `INH(p852) : f873;
        f873 = (f873 > p853) ? p853 : f873;
        f874 = 4095;
        f874 = (f874 >= `INH(p108)) ? `INH(p108) : f874;
        f874 = (f874 > p847) ? p847 : f874;
        f874 = (f874 > p851) ? p851 : f874;
        f875 = 4095;
        f875 = (f875 > p844) ? p844 : f875;
        f875 = (f875 >= `INH(p849)) ? `INH(p849) : f875;
        f875 = (f875 >= `INH(p853)) ? `INH(p853) : f875;
        f876 = 4095;
        f876 = (f876 > p843) ? p843 : f876;
        f876 = (f876 >= `INH(p854)) ? `INH(p854) : f876;
        f877 = 4095;
        f877 = (f877 > p120) ? p120 : f877;
        f877 = (f877 >= `INH(p845)) ? `INH(p845) : f877;
        f878 = 4095;
        f878 = (f878 >= `INH(p120)) ? `INH(p120) : f878;
        f878 = (f878 >= `INH(p845)) ? `INH(p845) : f878;
        f878 = (f878 > p854) ? p854 : f878;
        f879 = 4095;
        f879 = (f879 > p109) ? p109 : f879;
        f879 = (f879 >= `INH(p843)) ? `INH(p843) : f879;
        f879 = (f879 >= `INH(p854)) ? `INH(p854) : f879;
        f880 = 4095;
        f880 = (f880 >= `INH(p856)) ? `INH(p856) : f880;
        f880 = (f880 >= `INH(p857)) ? `INH(p857) : f880;
        f880 = (f880 > p861) ? p861 : f880;
        f881 = 4095;
        f881 = (f881 > p855) ? p855 : f881;
        f881 = (f881 >= `INH(p861)) ? `INH(p861) : f881;
        f882 = 4095;
        f882 = (f882 > p859) ? p859 : f882;
        f882 = (f882 >= `INH(p861)) ? `INH(p861) : f882;
        f883 = 4095;
        f883 = (f883 >= p856/2) ? p856/2 : f883;
        f883 = (f883 >= `INH(p860)) ? `INH(p860) : f883;
        f884 = 4095;
        f884 = (f884 >= `INH(p860)) ? `INH(p860) : f884;
        f884 = (f884 > p863) ? p863 : f884;
        f885 = 4095;
        f885 = (f885 > p856) ? p856 : f885;
        f885 = (f885 >= `INH(p863)) ? `INH(p863) : f885;
        f885 = (f885 > p865) ? p865 : f885;
        f886 = 4095;
        f886 = (f886 >= `INH(p863)) ? `INH(p863) : f886;
        f886 = (f886 > p866) ? p866 : f886;
        f887 = 4095;
        f887 = (f887 > p855) ? p855 : f887;
        f887 = (f887 >= `INH(p865)) ? `INH(p865) : f887;
        f887 = (f887 >= `INH(p866)) ? `INH(p866) : f887;
        f888 = 4095;
        f888 = (f888 > p855) ? p855 : f888;
        f888 = (f888 >= `INH(p864)) ? `INH(p864) : f888;
        f888 = (f888 >= `INH(p866)) ? `INH(p866) : f888;
        f889 = 4095;
        f889 = (f889 >= `INH(p866)) ? `INH(p866) : f889;
        f889 = (f889 > p868) ? p868 : f889;
        f890 = 4095;
        f890 = (f890 > p862) ? p862 : f890;
        f890 = (f890 >= `INH(p868)) ? `INH(p868) : f890;
        f891 = 4095;
        f891 = (f891 >= `INH(p868)) ? `INH(p868) : f891;
        f891 = (f891 > p869) ? p869 : f891;
        f892 = 4095;
        f892 = (f892 > p867) ? p867 : f892;
        f892 = (f892 >= `INH(p869)) ? `INH(p869) : f892;
        f893 = 4095;
        f893 = (f893 > p857) ? p857 : f893;
        f893 = (f893 > p864) ? p864 : f893;
        f893 = (f893 >= `INH(p865)) ? `INH(p865) : f893;
        f893 = (f893 >= `INH(p869)) ? `INH(p869) : f893;
        f894 = 4095;
        f894 = (f894 > p857) ? p857 : f894;
        f894 = (f894 >= `INH(p864)) ? `INH(p864) : f894;
        f894 = (f894 >= `INH(p869)) ? `INH(p869) : f894;
        f895 = 4095;
        f895 = (f895 > p127) ? p127 : f895;
        f895 = (f895 >= `INH(p871)) ? `INH(p871) : f895;
        f896 = 4095;
        f896 = (f896 > p870) ? p870 : f896;
        f896 = (f896 >= `INH(p872)) ? `INH(p872) : f896;
        f897 = 4095;
        f897 = (f897 >= `INH(p127)) ? `INH(p127) : f897;
        f897 = (f897 >= `INH(p871)) ? `INH(p871) : f897;
        f897 = (f897 > p872) ? p872 : f897;
        f898 = 4095;
        f898 = (f898 >= `INH(p870)) ? `INH(p870) : f898;
        f898 = (f898 >= `INH(p872)) ? `INH(p872) : f898;
        f898 = (f898 > p873) ? p873 : f898;
        f899 = 4095;
        f899 = (f899 > p128) ? p128 : f899;
        f899 = (f899 >= `INH(p875)) ? `INH(p875) : f899;
        f900 = 4095;
        f900 = (f900 > p874) ? p874 : f900;
        f900 = (f900 >= `INH(p876)) ? `INH(p876) : f900;
        f901 = 4095;
        f901 = (f901 >= `INH(p128)) ? `INH(p128) : f901;
        f901 = (f901 >= `INH(p875)) ? `INH(p875) : f901;
        f901 = (f901 > p876) ? p876 : f901;
        f902 = 4095;
        f902 = (f902 >= `INH(p874)) ? `INH(p874) : f902;
        f902 = (f902 >= `INH(p876)) ? `INH(p876) : f902;
        f902 = (f902 > p877) ? p877 : f902;
        f903 = 4095;
        f903 = (f903 >= `INH(p121)) ? `INH(p121) : f903;
        f903 = (f903 > p871) ? p871 : f903;
        f903 = (f903 > p875) ? p875 : f903;
        f904 = 4095;
        f904 = (f904 > p857) ? p857 : f904;
        f904 = (f904 >= `INH(p873)) ? `INH(p873) : f904;
        f904 = (f904 >= `INH(p877)) ? `INH(p877) : f904;
        f905 = 4095;
        f905 = (f905 > p858) ? p858 : f905;
        f905 = (f905 >= `INH(p878)) ? `INH(p878) : f905;
        f906 = 4095;
        f906 = (f906 > p129) ? p129 : f906;
        f906 = (f906 >= `INH(p859)) ? `INH(p859) : f906;
        f907 = 4095;
        f907 = (f907 >= `INH(p129)) ? `INH(p129) : f907;
        f907 = (f907 >= `INH(p859)) ? `INH(p859) : f907;
        f907 = (f907 > p878) ? p878 : f907;
        f908 = 4095;
        f908 = (f908 > p122) ? p122 : f908;
        f908 = (f908 >= `INH(p858)) ? `INH(p858) : f908;
        f908 = (f908 >= `INH(p878)) ? `INH(p878) : f908;
        f909 = 4095;
        f909 = (f909 >= `INH(p880)) ? `INH(p880) : f909;
        f909 = (f909 >= `INH(p881)) ? `INH(p881) : f909;
        f909 = (f909 > p885) ? p885 : f909;
        f910 = 4095;
        f910 = (f910 > p879) ? p879 : f910;
        f910 = (f910 >= `INH(p885)) ? `INH(p885) : f910;
        f911 = 4095;
        f911 = (f911 > p883) ? p883 : f911;
        f911 = (f911 >= `INH(p885)) ? `INH(p885) : f911;
        f912 = 4095;
        f912 = (f912 >= p880/2) ? p880/2 : f912;
        f912 = (f912 >= `INH(p884)) ? `INH(p884) : f912;
        f913 = 4095;
        f913 = (f913 >= `INH(p884)) ? `INH(p884) : f913;
        f913 = (f913 > p887) ? p887 : f913;
        f914 = 4095;
        f914 = (f914 > p880) ? p880 : f914;
        f914 = (f914 >= `INH(p887)) ? `INH(p887) : f914;
        f914 = (f914 > p889) ? p889 : f914;
        f915 = 4095;
        f915 = (f915 >= `INH(p887)) ? `INH(p887) : f915;
        f915 = (f915 > p890) ? p890 : f915;
        f916 = 4095;
        f916 = (f916 > p879) ? p879 : f916;
        f916 = (f916 >= `INH(p889)) ? `INH(p889) : f916;
        f916 = (f916 >= `INH(p890)) ? `INH(p890) : f916;
        f917 = 4095;
        f917 = (f917 > p879) ? p879 : f917;
        f917 = (f917 >= `INH(p888)) ? `INH(p888) : f917;
        f917 = (f917 >= `INH(p890)) ? `INH(p890) : f917;
        f918 = 4095;
        f918 = (f918 >= `INH(p890)) ? `INH(p890) : f918;
        f918 = (f918 > p892) ? p892 : f918;
        f919 = 4095;
        f919 = (f919 > p886) ? p886 : f919;
        f919 = (f919 >= `INH(p892)) ? `INH(p892) : f919;
        f920 = 4095;
        f920 = (f920 >= `INH(p892)) ? `INH(p892) : f920;
        f920 = (f920 > p893) ? p893 : f920;
        f921 = 4095;
        f921 = (f921 > p891) ? p891 : f921;
        f921 = (f921 >= `INH(p893)) ? `INH(p893) : f921;
        f922 = 4095;
        f922 = (f922 > p881) ? p881 : f922;
        f922 = (f922 > p888) ? p888 : f922;
        f922 = (f922 >= `INH(p889)) ? `INH(p889) : f922;
        f922 = (f922 >= `INH(p893)) ? `INH(p893) : f922;
        f923 = 4095;
        f923 = (f923 > p881) ? p881 : f923;
        f923 = (f923 >= `INH(p888)) ? `INH(p888) : f923;
        f923 = (f923 >= `INH(p893)) ? `INH(p893) : f923;
        f924 = 4095;
        f924 = (f924 > p130) ? p130 : f924;
        f924 = (f924 >= `INH(p895)) ? `INH(p895) : f924;
        f925 = 4095;
        f925 = (f925 > p894) ? p894 : f925;
        f925 = (f925 >= `INH(p896)) ? `INH(p896) : f925;
        f926 = 4095;
        f926 = (f926 >= `INH(p130)) ? `INH(p130) : f926;
        f926 = (f926 >= `INH(p895)) ? `INH(p895) : f926;
        f926 = (f926 > p896) ? p896 : f926;
        f927 = 4095;
        f927 = (f927 >= `INH(p894)) ? `INH(p894) : f927;
        f927 = (f927 >= `INH(p896)) ? `INH(p896) : f927;
        f927 = (f927 > p897) ? p897 : f927;
        f928 = 4095;
        f928 = (f928 > p131) ? p131 : f928;
        f928 = (f928 >= `INH(p899)) ? `INH(p899) : f928;
        f929 = 4095;
        f929 = (f929 > p898) ? p898 : f929;
        f929 = (f929 >= `INH(p900)) ? `INH(p900) : f929;
        f930 = 4095;
        f930 = (f930 >= `INH(p131)) ? `INH(p131) : f930;
        f930 = (f930 >= `INH(p899)) ? `INH(p899) : f930;
        f930 = (f930 > p900) ? p900 : f930;
        f931 = 4095;
        f931 = (f931 >= `INH(p898)) ? `INH(p898) : f931;
        f931 = (f931 >= `INH(p900)) ? `INH(p900) : f931;
        f931 = (f931 > p901) ? p901 : f931;
        f932 = 4095;
        f932 = (f932 >= `INH(p122)) ? `INH(p122) : f932;
        f932 = (f932 > p895) ? p895 : f932;
        f932 = (f932 > p899) ? p899 : f932;
        f933 = 4095;
        f933 = (f933 > p881) ? p881 : f933;
        f933 = (f933 >= `INH(p897)) ? `INH(p897) : f933;
        f933 = (f933 >= `INH(p901)) ? `INH(p901) : f933;
        f934 = 4095;
        f934 = (f934 > p882) ? p882 : f934;
        f934 = (f934 >= `INH(p902)) ? `INH(p902) : f934;
        f935 = 4095;
        f935 = (f935 > p132) ? p132 : f935;
        f935 = (f935 >= `INH(p883)) ? `INH(p883) : f935;
        f936 = 4095;
        f936 = (f936 >= `INH(p132)) ? `INH(p132) : f936;
        f936 = (f936 >= `INH(p883)) ? `INH(p883) : f936;
        f936 = (f936 > p902) ? p902 : f936;
        f937 = 4095;
        f937 = (f937 > p123) ? p123 : f937;
        f937 = (f937 >= `INH(p882)) ? `INH(p882) : f937;
        f937 = (f937 >= `INH(p902)) ? `INH(p902) : f937;
        f938 = 4095;
        f938 = (f938 > p904) ? p904 : f938;
        f938 = (f938 >= `INH(p906)) ? `INH(p906) : f938;
        f939 = 4095;
        f939 = (f939 >= `INH(p903)) ? `INH(p903) : f939;
        f939 = (f939 >= `INH(p904)) ? `INH(p904) : f939;
        f939 = (f939 >= `INH(p906)) ? `INH(p906) : f939;
        f939 = (f939 > p907) ? p907 : f939;
        f940 = 4095;
        f940 = (f940 > p129) ? p129 : f940;
        f940 = (f940 >= `INH(p909)) ? `INH(p909) : f940;
        f941 = 4095;
        f941 = (f941 > p908) ? p908 : f941;
        f941 = (f941 >= `INH(p910)) ? `INH(p910) : f941;
        f942 = 4095;
        f942 = (f942 >= `INH(p129)) ? `INH(p129) : f942;
        f942 = (f942 >= `INH(p909)) ? `INH(p909) : f942;
        f942 = (f942 > p910) ? p910 : f942;
        f943 = 4095;
        f943 = (f943 >= `INH(p908)) ? `INH(p908) : f943;
        f943 = (f943 >= `INH(p910)) ? `INH(p910) : f943;
        f943 = (f943 > p911) ? p911 : f943;
        f944 = 4095;
        f944 = (f944 > p132) ? p132 : f944;
        f944 = (f944 >= `INH(p913)) ? `INH(p913) : f944;
        f945 = 4095;
        f945 = (f945 > p912) ? p912 : f945;
        f945 = (f945 >= `INH(p914)) ? `INH(p914) : f945;
        f946 = 4095;
        f946 = (f946 >= `INH(p132)) ? `INH(p132) : f946;
        f946 = (f946 >= `INH(p913)) ? `INH(p913) : f946;
        f946 = (f946 > p914) ? p914 : f946;
        f947 = 4095;
        f947 = (f947 >= `INH(p912)) ? `INH(p912) : f947;
        f947 = (f947 >= `INH(p914)) ? `INH(p914) : f947;
        f947 = (f947 > p915) ? p915 : f947;
        f948 = 4095;
        f948 = (f948 >= `INH(p123)) ? `INH(p123) : f948;
        f948 = (f948 > p909) ? p909 : f948;
        f948 = (f948 > p913) ? p913 : f948;
        f949 = 4095;
        f949 = (f949 > p906) ? p906 : f949;
        f949 = (f949 >= `INH(p911)) ? `INH(p911) : f949;
        f949 = (f949 >= `INH(p915)) ? `INH(p915) : f949;
        f950 = 4095;
        f950 = (f950 > p905) ? p905 : f950;
        f950 = (f950 >= `INH(p916)) ? `INH(p916) : f950;
        f951 = 4095;
        f951 = (f951 > p133) ? p133 : f951;
        f951 = (f951 >= `INH(p907)) ? `INH(p907) : f951;
        f952 = 4095;
        f952 = (f952 >= `INH(p133)) ? `INH(p133) : f952;
        f952 = (f952 >= `INH(p907)) ? `INH(p907) : f952;
        f952 = (f952 > p916) ? p916 : f952;
        f953 = 4095;
        f953 = (f953 > p124) ? p124 : f953;
        f953 = (f953 >= `INH(p905)) ? `INH(p905) : f953;
        f953 = (f953 >= `INH(p916)) ? `INH(p916) : f953;
        f954 = 4095;
        f954 = (f954 >= `INH(p918)) ? `INH(p918) : f954;
        f954 = (f954 >= `INH(p919)) ? `INH(p919) : f954;
        f954 = (f954 > p923) ? p923 : f954;
        f955 = 4095;
        f955 = (f955 > p917) ? p917 : f955;
        f955 = (f955 >= `INH(p923)) ? `INH(p923) : f955;
        f956 = 4095;
        f956 = (f956 > p921) ? p921 : f956;
        f956 = (f956 >= `INH(p923)) ? `INH(p923) : f956;
        f957 = 4095;
        f957 = (f957 >= p918/2) ? p918/2 : f957;
        f957 = (f957 >= `INH(p922)) ? `INH(p922) : f957;
        f958 = 4095;
        f958 = (f958 >= `INH(p922)) ? `INH(p922) : f958;
        f958 = (f958 > p925) ? p925 : f958;
        f959 = 4095;
        f959 = (f959 > p918) ? p918 : f959;
        f959 = (f959 >= `INH(p925)) ? `INH(p925) : f959;
        f959 = (f959 > p927) ? p927 : f959;
        f960 = 4095;
        f960 = (f960 >= `INH(p925)) ? `INH(p925) : f960;
        f960 = (f960 > p928) ? p928 : f960;
        f961 = 4095;
        f961 = (f961 > p917) ? p917 : f961;
        f961 = (f961 >= `INH(p927)) ? `INH(p927) : f961;
        f961 = (f961 >= `INH(p928)) ? `INH(p928) : f961;
        f962 = 4095;
        f962 = (f962 > p917) ? p917 : f962;
        f962 = (f962 >= `INH(p926)) ? `INH(p926) : f962;
        f962 = (f962 >= `INH(p928)) ? `INH(p928) : f962;
        f963 = 4095;
        f963 = (f963 >= `INH(p928)) ? `INH(p928) : f963;
        f963 = (f963 > p930) ? p930 : f963;
        f964 = 4095;
        f964 = (f964 > p924) ? p924 : f964;
        f964 = (f964 >= `INH(p930)) ? `INH(p930) : f964;
        f965 = 4095;
        f965 = (f965 >= `INH(p930)) ? `INH(p930) : f965;
        f965 = (f965 > p931) ? p931 : f965;
        f966 = 4095;
        f966 = (f966 > p929) ? p929 : f966;
        f966 = (f966 >= `INH(p931)) ? `INH(p931) : f966;
        f967 = 4095;
        f967 = (f967 > p919) ? p919 : f967;
        f967 = (f967 > p926) ? p926 : f967;
        f967 = (f967 >= `INH(p927)) ? `INH(p927) : f967;
        f967 = (f967 >= `INH(p931)) ? `INH(p931) : f967;
        f968 = 4095;
        f968 = (f968 > p919) ? p919 : f968;
        f968 = (f968 >= `INH(p926)) ? `INH(p926) : f968;
        f968 = (f968 >= `INH(p931)) ? `INH(p931) : f968;
        f969 = 4095;
        f969 = (f969 > p134) ? p134 : f969;
        f969 = (f969 >= `INH(p933)) ? `INH(p933) : f969;
        f970 = 4095;
        f970 = (f970 > p932) ? p932 : f970;
        f970 = (f970 >= `INH(p934)) ? `INH(p934) : f970;
        f971 = 4095;
        f971 = (f971 >= `INH(p134)) ? `INH(p134) : f971;
        f971 = (f971 >= `INH(p933)) ? `INH(p933) : f971;
        f971 = (f971 > p934) ? p934 : f971;
        f972 = 4095;
        f972 = (f972 >= `INH(p932)) ? `INH(p932) : f972;
        f972 = (f972 >= `INH(p934)) ? `INH(p934) : f972;
        f972 = (f972 > p935) ? p935 : f972;
        f973 = 4095;
        f973 = (f973 > p135) ? p135 : f973;
        f973 = (f973 >= `INH(p937)) ? `INH(p937) : f973;
        f974 = 4095;
        f974 = (f974 > p936) ? p936 : f974;
        f974 = (f974 >= `INH(p938)) ? `INH(p938) : f974;
        f975 = 4095;
        f975 = (f975 >= `INH(p135)) ? `INH(p135) : f975;
        f975 = (f975 >= `INH(p937)) ? `INH(p937) : f975;
        f975 = (f975 > p938) ? p938 : f975;
        f976 = 4095;
        f976 = (f976 >= `INH(p936)) ? `INH(p936) : f976;
        f976 = (f976 >= `INH(p938)) ? `INH(p938) : f976;
        f976 = (f976 > p939) ? p939 : f976;
        f977 = 4095;
        f977 = (f977 >= `INH(p124)) ? `INH(p124) : f977;
        f977 = (f977 > p933) ? p933 : f977;
        f977 = (f977 > p937) ? p937 : f977;
        f978 = 4095;
        f978 = (f978 > p919) ? p919 : f978;
        f978 = (f978 >= `INH(p935)) ? `INH(p935) : f978;
        f978 = (f978 >= `INH(p939)) ? `INH(p939) : f978;
        f979 = 4095;
        f979 = (f979 > p920) ? p920 : f979;
        f979 = (f979 >= `INH(p940)) ? `INH(p940) : f979;
        f980 = 4095;
        f980 = (f980 > p136) ? p136 : f980;
        f980 = (f980 >= `INH(p921)) ? `INH(p921) : f980;
        f981 = 4095;
        f981 = (f981 >= `INH(p136)) ? `INH(p136) : f981;
        f981 = (f981 >= `INH(p921)) ? `INH(p921) : f981;
        f981 = (f981 > p940) ? p940 : f981;
        f982 = 4095;
        f982 = (f982 > p125) ? p125 : f982;
        f982 = (f982 >= `INH(p920)) ? `INH(p920) : f982;
        f982 = (f982 >= `INH(p940)) ? `INH(p940) : f982;
        f983 = 4095;
        f983 = (f983 > p942) ? p942 : f983;
        f983 = (f983 >= `INH(p944)) ? `INH(p944) : f983;
        f984 = 4095;
        f984 = (f984 >= `INH(p941)) ? `INH(p941) : f984;
        f984 = (f984 >= `INH(p942)) ? `INH(p942) : f984;
        f984 = (f984 >= `INH(p944)) ? `INH(p944) : f984;
        f984 = (f984 > p945) ? p945 : f984;
        f985 = 4095;
        f985 = (f985 > p133) ? p133 : f985;
        f985 = (f985 >= `INH(p947)) ? `INH(p947) : f985;
        f986 = 4095;
        f986 = (f986 > p946) ? p946 : f986;
        f986 = (f986 >= `INH(p948)) ? `INH(p948) : f986;
        f987 = 4095;
        f987 = (f987 >= `INH(p133)) ? `INH(p133) : f987;
        f987 = (f987 >= `INH(p947)) ? `INH(p947) : f987;
        f987 = (f987 > p948) ? p948 : f987;
        f988 = 4095;
        f988 = (f988 >= `INH(p946)) ? `INH(p946) : f988;
        f988 = (f988 >= `INH(p948)) ? `INH(p948) : f988;
        f988 = (f988 > p949) ? p949 : f988;
        f989 = 4095;
        f989 = (f989 > p136) ? p136 : f989;
        f989 = (f989 >= `INH(p951)) ? `INH(p951) : f989;
        f990 = 4095;
        f990 = (f990 > p950) ? p950 : f990;
        f990 = (f990 >= `INH(p952)) ? `INH(p952) : f990;
        f991 = 4095;
        f991 = (f991 >= `INH(p136)) ? `INH(p136) : f991;
        f991 = (f991 >= `INH(p951)) ? `INH(p951) : f991;
        f991 = (f991 > p952) ? p952 : f991;
        f992 = 4095;
        f992 = (f992 >= `INH(p950)) ? `INH(p950) : f992;
        f992 = (f992 >= `INH(p952)) ? `INH(p952) : f992;
        f992 = (f992 > p953) ? p953 : f992;
        f993 = 4095;
        f993 = (f993 >= `INH(p125)) ? `INH(p125) : f993;
        f993 = (f993 > p947) ? p947 : f993;
        f993 = (f993 > p951) ? p951 : f993;
        f994 = 4095;
        f994 = (f994 > p944) ? p944 : f994;
        f994 = (f994 >= `INH(p949)) ? `INH(p949) : f994;
        f994 = (f994 >= `INH(p953)) ? `INH(p953) : f994;
        f995 = 4095;
        f995 = (f995 > p943) ? p943 : f995;
        f995 = (f995 >= `INH(p954)) ? `INH(p954) : f995;
        f996 = 4095;
        f996 = (f996 > p137) ? p137 : f996;
        f996 = (f996 >= `INH(p945)) ? `INH(p945) : f996;
        f997 = 4095;
        f997 = (f997 >= `INH(p137)) ? `INH(p137) : f997;
        f997 = (f997 >= `INH(p945)) ? `INH(p945) : f997;
        f997 = (f997 > p954) ? p954 : f997;
        f998 = 4095;
        f998 = (f998 > p126) ? p126 : f998;
        f998 = (f998 >= `INH(p943)) ? `INH(p943) : f998;
        f998 = (f998 >= `INH(p954)) ? `INH(p954) : f998;
        f999 = 4095;
        f999 = (f999 >= `INH(p956)) ? `INH(p956) : f999;
        f999 = (f999 >= `INH(p957)) ? `INH(p957) : f999;
        f999 = (f999 > p961) ? p961 : f999;
        f1000 = 4095;
        f1000 = (f1000 > p955) ? p955 : f1000;
        f1000 = (f1000 >= `INH(p961)) ? `INH(p961) : f1000;
        f1001 = 4095;
        f1001 = (f1001 > p959) ? p959 : f1001;
        f1001 = (f1001 >= `INH(p961)) ? `INH(p961) : f1001;
        f1002 = 4095;
        f1002 = (f1002 >= p956/2) ? p956/2 : f1002;
        f1002 = (f1002 >= `INH(p960)) ? `INH(p960) : f1002;
        f1003 = 4095;
        f1003 = (f1003 >= `INH(p960)) ? `INH(p960) : f1003;
        f1003 = (f1003 > p963) ? p963 : f1003;
        f1004 = 4095;
        f1004 = (f1004 > p956) ? p956 : f1004;
        f1004 = (f1004 >= `INH(p963)) ? `INH(p963) : f1004;
        f1004 = (f1004 > p965) ? p965 : f1004;
        f1005 = 4095;
        f1005 = (f1005 >= `INH(p963)) ? `INH(p963) : f1005;
        f1005 = (f1005 > p966) ? p966 : f1005;
        f1006 = 4095;
        f1006 = (f1006 > p955) ? p955 : f1006;
        f1006 = (f1006 >= `INH(p965)) ? `INH(p965) : f1006;
        f1006 = (f1006 >= `INH(p966)) ? `INH(p966) : f1006;
        f1007 = 4095;
        f1007 = (f1007 > p955) ? p955 : f1007;
        f1007 = (f1007 >= `INH(p964)) ? `INH(p964) : f1007;
        f1007 = (f1007 >= `INH(p966)) ? `INH(p966) : f1007;
        f1008 = 4095;
        f1008 = (f1008 >= `INH(p966)) ? `INH(p966) : f1008;
        f1008 = (f1008 > p968) ? p968 : f1008;
        f1009 = 4095;
        f1009 = (f1009 > p962) ? p962 : f1009;
        f1009 = (f1009 >= `INH(p968)) ? `INH(p968) : f1009;
        f1010 = 4095;
        f1010 = (f1010 >= `INH(p968)) ? `INH(p968) : f1010;
        f1010 = (f1010 > p969) ? p969 : f1010;
        f1011 = 4095;
        f1011 = (f1011 > p967) ? p967 : f1011;
        f1011 = (f1011 >= `INH(p969)) ? `INH(p969) : f1011;
        f1012 = 4095;
        f1012 = (f1012 > p957) ? p957 : f1012;
        f1012 = (f1012 > p964) ? p964 : f1012;
        f1012 = (f1012 >= `INH(p965)) ? `INH(p965) : f1012;
        f1012 = (f1012 >= `INH(p969)) ? `INH(p969) : f1012;
        f1013 = 4095;
        f1013 = (f1013 > p957) ? p957 : f1013;
        f1013 = (f1013 >= `INH(p964)) ? `INH(p964) : f1013;
        f1013 = (f1013 >= `INH(p969)) ? `INH(p969) : f1013;
        f1014 = 4095;
        f1014 = (f1014 > p144) ? p144 : f1014;
        f1014 = (f1014 >= `INH(p971)) ? `INH(p971) : f1014;
        f1015 = 4095;
        f1015 = (f1015 > p970) ? p970 : f1015;
        f1015 = (f1015 >= `INH(p972)) ? `INH(p972) : f1015;
        f1016 = 4095;
        f1016 = (f1016 >= `INH(p144)) ? `INH(p144) : f1016;
        f1016 = (f1016 >= `INH(p971)) ? `INH(p971) : f1016;
        f1016 = (f1016 > p972) ? p972 : f1016;
        f1017 = 4095;
        f1017 = (f1017 >= `INH(p970)) ? `INH(p970) : f1017;
        f1017 = (f1017 >= `INH(p972)) ? `INH(p972) : f1017;
        f1017 = (f1017 > p973) ? p973 : f1017;
        f1018 = 4095;
        f1018 = (f1018 > p145) ? p145 : f1018;
        f1018 = (f1018 >= `INH(p975)) ? `INH(p975) : f1018;
        f1019 = 4095;
        f1019 = (f1019 > p974) ? p974 : f1019;
        f1019 = (f1019 >= `INH(p976)) ? `INH(p976) : f1019;
        f1020 = 4095;
        f1020 = (f1020 >= `INH(p145)) ? `INH(p145) : f1020;
        f1020 = (f1020 >= `INH(p975)) ? `INH(p975) : f1020;
        f1020 = (f1020 > p976) ? p976 : f1020;
        f1021 = 4095;
        f1021 = (f1021 >= `INH(p974)) ? `INH(p974) : f1021;
        f1021 = (f1021 >= `INH(p976)) ? `INH(p976) : f1021;
        f1021 = (f1021 > p977) ? p977 : f1021;
        f1022 = 4095;
        f1022 = (f1022 >= `INH(p138)) ? `INH(p138) : f1022;
        f1022 = (f1022 > p971) ? p971 : f1022;
        f1022 = (f1022 > p975) ? p975 : f1022;
        f1023 = 4095;
        f1023 = (f1023 > p957) ? p957 : f1023;
        f1023 = (f1023 >= `INH(p973)) ? `INH(p973) : f1023;
        f1023 = (f1023 >= `INH(p977)) ? `INH(p977) : f1023;
        f1024 = 4095;
        f1024 = (f1024 > p958) ? p958 : f1024;
        f1024 = (f1024 >= `INH(p978)) ? `INH(p978) : f1024;
        f1025 = 4095;
        f1025 = (f1025 > p146) ? p146 : f1025;
        f1025 = (f1025 >= `INH(p959)) ? `INH(p959) : f1025;
        f1026 = 4095;
        f1026 = (f1026 >= `INH(p146)) ? `INH(p146) : f1026;
        f1026 = (f1026 >= `INH(p959)) ? `INH(p959) : f1026;
        f1026 = (f1026 > p978) ? p978 : f1026;
        f1027 = 4095;
        f1027 = (f1027 > p139) ? p139 : f1027;
        f1027 = (f1027 >= `INH(p958)) ? `INH(p958) : f1027;
        f1027 = (f1027 >= `INH(p978)) ? `INH(p978) : f1027;
        f1028 = 4095;
        f1028 = (f1028 >= `INH(p980)) ? `INH(p980) : f1028;
        f1028 = (f1028 >= `INH(p981)) ? `INH(p981) : f1028;
        f1028 = (f1028 > p985) ? p985 : f1028;
        f1029 = 4095;
        f1029 = (f1029 > p979) ? p979 : f1029;
        f1029 = (f1029 >= `INH(p985)) ? `INH(p985) : f1029;
        f1030 = 4095;
        f1030 = (f1030 > p983) ? p983 : f1030;
        f1030 = (f1030 >= `INH(p985)) ? `INH(p985) : f1030;
        f1031 = 4095;
        f1031 = (f1031 >= p980/2) ? p980/2 : f1031;
        f1031 = (f1031 >= `INH(p984)) ? `INH(p984) : f1031;
        f1032 = 4095;
        f1032 = (f1032 >= `INH(p984)) ? `INH(p984) : f1032;
        f1032 = (f1032 > p987) ? p987 : f1032;
        f1033 = 4095;
        f1033 = (f1033 > p980) ? p980 : f1033;
        f1033 = (f1033 >= `INH(p987)) ? `INH(p987) : f1033;
        f1033 = (f1033 > p989) ? p989 : f1033;
        f1034 = 4095;
        f1034 = (f1034 >= `INH(p987)) ? `INH(p987) : f1034;
        f1034 = (f1034 > p990) ? p990 : f1034;
        f1035 = 4095;
        f1035 = (f1035 > p979) ? p979 : f1035;
        f1035 = (f1035 >= `INH(p989)) ? `INH(p989) : f1035;
        f1035 = (f1035 >= `INH(p990)) ? `INH(p990) : f1035;
        f1036 = 4095;
        f1036 = (f1036 > p979) ? p979 : f1036;
        f1036 = (f1036 >= `INH(p988)) ? `INH(p988) : f1036;
        f1036 = (f1036 >= `INH(p990)) ? `INH(p990) : f1036;
        f1037 = 4095;
        f1037 = (f1037 >= `INH(p990)) ? `INH(p990) : f1037;
        f1037 = (f1037 > p992) ? p992 : f1037;
        f1038 = 4095;
        f1038 = (f1038 > p986) ? p986 : f1038;
        f1038 = (f1038 >= `INH(p992)) ? `INH(p992) : f1038;
        f1039 = 4095;
        f1039 = (f1039 >= `INH(p992)) ? `INH(p992) : f1039;
        f1039 = (f1039 > p993) ? p993 : f1039;
        f1040 = 4095;
        f1040 = (f1040 > p991) ? p991 : f1040;
        f1040 = (f1040 >= `INH(p993)) ? `INH(p993) : f1040;
        f1041 = 4095;
        f1041 = (f1041 > p981) ? p981 : f1041;
        f1041 = (f1041 > p988) ? p988 : f1041;
        f1041 = (f1041 >= `INH(p989)) ? `INH(p989) : f1041;
        f1041 = (f1041 >= `INH(p993)) ? `INH(p993) : f1041;
        f1042 = 4095;
        f1042 = (f1042 > p981) ? p981 : f1042;
        f1042 = (f1042 >= `INH(p988)) ? `INH(p988) : f1042;
        f1042 = (f1042 >= `INH(p993)) ? `INH(p993) : f1042;
        f1043 = 4095;
        f1043 = (f1043 > p147) ? p147 : f1043;
        f1043 = (f1043 >= `INH(p995)) ? `INH(p995) : f1043;
        f1044 = 4095;
        f1044 = (f1044 > p994) ? p994 : f1044;
        f1044 = (f1044 >= `INH(p996)) ? `INH(p996) : f1044;
        f1045 = 4095;
        f1045 = (f1045 >= `INH(p147)) ? `INH(p147) : f1045;
        f1045 = (f1045 >= `INH(p995)) ? `INH(p995) : f1045;
        f1045 = (f1045 > p996) ? p996 : f1045;
        f1046 = 4095;
        f1046 = (f1046 >= `INH(p994)) ? `INH(p994) : f1046;
        f1046 = (f1046 >= `INH(p996)) ? `INH(p996) : f1046;
        f1046 = (f1046 > p997) ? p997 : f1046;
        f1047 = 4095;
        f1047 = (f1047 > p148) ? p148 : f1047;
        f1047 = (f1047 >= `INH(p999)) ? `INH(p999) : f1047;
        f1048 = 4095;
        f1048 = (f1048 > p998) ? p998 : f1048;
        f1048 = (f1048 >= `INH(p1000)) ? `INH(p1000) : f1048;
        f1049 = 4095;
        f1049 = (f1049 >= `INH(p148)) ? `INH(p148) : f1049;
        f1049 = (f1049 >= `INH(p999)) ? `INH(p999) : f1049;
        f1049 = (f1049 > p1000) ? p1000 : f1049;
        f1050 = 4095;
        f1050 = (f1050 >= `INH(p998)) ? `INH(p998) : f1050;
        f1050 = (f1050 >= `INH(p1000)) ? `INH(p1000) : f1050;
        f1050 = (f1050 > p1001) ? p1001 : f1050;
        f1051 = 4095;
        f1051 = (f1051 >= `INH(p139)) ? `INH(p139) : f1051;
        f1051 = (f1051 > p995) ? p995 : f1051;
        f1051 = (f1051 > p999) ? p999 : f1051;
        f1052 = 4095;
        f1052 = (f1052 > p981) ? p981 : f1052;
        f1052 = (f1052 >= `INH(p997)) ? `INH(p997) : f1052;
        f1052 = (f1052 >= `INH(p1001)) ? `INH(p1001) : f1052;
        f1053 = 4095;
        f1053 = (f1053 > p982) ? p982 : f1053;
        f1053 = (f1053 >= `INH(p1002)) ? `INH(p1002) : f1053;
        f1054 = 4095;
        f1054 = (f1054 > p149) ? p149 : f1054;
        f1054 = (f1054 >= `INH(p983)) ? `INH(p983) : f1054;
        f1055 = 4095;
        f1055 = (f1055 >= `INH(p149)) ? `INH(p149) : f1055;
        f1055 = (f1055 >= `INH(p983)) ? `INH(p983) : f1055;
        f1055 = (f1055 > p1002) ? p1002 : f1055;
        f1056 = 4095;
        f1056 = (f1056 > p140) ? p140 : f1056;
        f1056 = (f1056 >= `INH(p982)) ? `INH(p982) : f1056;
        f1056 = (f1056 >= `INH(p1002)) ? `INH(p1002) : f1056;
        f1057 = 4095;
        f1057 = (f1057 > p1004) ? p1004 : f1057;
        f1057 = (f1057 >= `INH(p1006)) ? `INH(p1006) : f1057;
        f1058 = 4095;
        f1058 = (f1058 >= `INH(p1003)) ? `INH(p1003) : f1058;
        f1058 = (f1058 >= `INH(p1004)) ? `INH(p1004) : f1058;
        f1058 = (f1058 >= `INH(p1006)) ? `INH(p1006) : f1058;
        f1058 = (f1058 > p1007) ? p1007 : f1058;
        f1059 = 4095;
        f1059 = (f1059 > p146) ? p146 : f1059;
        f1059 = (f1059 >= `INH(p1009)) ? `INH(p1009) : f1059;
        f1060 = 4095;
        f1060 = (f1060 > p1008) ? p1008 : f1060;
        f1060 = (f1060 >= `INH(p1010)) ? `INH(p1010) : f1060;
        f1061 = 4095;
        f1061 = (f1061 >= `INH(p146)) ? `INH(p146) : f1061;
        f1061 = (f1061 >= `INH(p1009)) ? `INH(p1009) : f1061;
        f1061 = (f1061 > p1010) ? p1010 : f1061;
        f1062 = 4095;
        f1062 = (f1062 >= `INH(p1008)) ? `INH(p1008) : f1062;
        f1062 = (f1062 >= `INH(p1010)) ? `INH(p1010) : f1062;
        f1062 = (f1062 > p1011) ? p1011 : f1062;
        f1063 = 4095;
        f1063 = (f1063 > p149) ? p149 : f1063;
        f1063 = (f1063 >= `INH(p1013)) ? `INH(p1013) : f1063;
        f1064 = 4095;
        f1064 = (f1064 > p1012) ? p1012 : f1064;
        f1064 = (f1064 >= `INH(p1014)) ? `INH(p1014) : f1064;
        f1065 = 4095;
        f1065 = (f1065 >= `INH(p149)) ? `INH(p149) : f1065;
        f1065 = (f1065 >= `INH(p1013)) ? `INH(p1013) : f1065;
        f1065 = (f1065 > p1014) ? p1014 : f1065;
        f1066 = 4095;
        f1066 = (f1066 >= `INH(p1012)) ? `INH(p1012) : f1066;
        f1066 = (f1066 >= `INH(p1014)) ? `INH(p1014) : f1066;
        f1066 = (f1066 > p1015) ? p1015 : f1066;
        f1067 = 4095;
        f1067 = (f1067 >= `INH(p140)) ? `INH(p140) : f1067;
        f1067 = (f1067 > p1009) ? p1009 : f1067;
        f1067 = (f1067 > p1013) ? p1013 : f1067;
        f1068 = 4095;
        f1068 = (f1068 > p1006) ? p1006 : f1068;
        f1068 = (f1068 >= `INH(p1011)) ? `INH(p1011) : f1068;
        f1068 = (f1068 >= `INH(p1015)) ? `INH(p1015) : f1068;
        f1069 = 4095;
        f1069 = (f1069 > p1005) ? p1005 : f1069;
        f1069 = (f1069 >= `INH(p1016)) ? `INH(p1016) : f1069;
        f1070 = 4095;
        f1070 = (f1070 > p150) ? p150 : f1070;
        f1070 = (f1070 >= `INH(p1007)) ? `INH(p1007) : f1070;
        f1071 = 4095;
        f1071 = (f1071 >= `INH(p150)) ? `INH(p150) : f1071;
        f1071 = (f1071 >= `INH(p1007)) ? `INH(p1007) : f1071;
        f1071 = (f1071 > p1016) ? p1016 : f1071;
        f1072 = 4095;
        f1072 = (f1072 > p141) ? p141 : f1072;
        f1072 = (f1072 >= `INH(p1005)) ? `INH(p1005) : f1072;
        f1072 = (f1072 >= `INH(p1016)) ? `INH(p1016) : f1072;
        f1073 = 4095;
        f1073 = (f1073 >= `INH(p1018)) ? `INH(p1018) : f1073;
        f1073 = (f1073 >= `INH(p1019)) ? `INH(p1019) : f1073;
        f1073 = (f1073 > p1023) ? p1023 : f1073;
        f1074 = 4095;
        f1074 = (f1074 > p1017) ? p1017 : f1074;
        f1074 = (f1074 >= `INH(p1023)) ? `INH(p1023) : f1074;
        f1075 = 4095;
        f1075 = (f1075 > p1021) ? p1021 : f1075;
        f1075 = (f1075 >= `INH(p1023)) ? `INH(p1023) : f1075;
        f1076 = 4095;
        f1076 = (f1076 >= p1018/2) ? p1018/2 : f1076;
        f1076 = (f1076 >= `INH(p1022)) ? `INH(p1022) : f1076;
        f1077 = 4095;
        f1077 = (f1077 >= `INH(p1022)) ? `INH(p1022) : f1077;
        f1077 = (f1077 > p1025) ? p1025 : f1077;
        f1078 = 4095;
        f1078 = (f1078 > p1018) ? p1018 : f1078;
        f1078 = (f1078 >= `INH(p1025)) ? `INH(p1025) : f1078;
        f1078 = (f1078 > p1027) ? p1027 : f1078;
        f1079 = 4095;
        f1079 = (f1079 >= `INH(p1025)) ? `INH(p1025) : f1079;
        f1079 = (f1079 > p1028) ? p1028 : f1079;
        f1080 = 4095;
        f1080 = (f1080 > p1017) ? p1017 : f1080;
        f1080 = (f1080 >= `INH(p1027)) ? `INH(p1027) : f1080;
        f1080 = (f1080 >= `INH(p1028)) ? `INH(p1028) : f1080;
        f1081 = 4095;
        f1081 = (f1081 > p1017) ? p1017 : f1081;
        f1081 = (f1081 >= `INH(p1026)) ? `INH(p1026) : f1081;
        f1081 = (f1081 >= `INH(p1028)) ? `INH(p1028) : f1081;
        f1082 = 4095;
        f1082 = (f1082 >= `INH(p1028)) ? `INH(p1028) : f1082;
        f1082 = (f1082 > p1030) ? p1030 : f1082;
        f1083 = 4095;
        f1083 = (f1083 > p1024) ? p1024 : f1083;
        f1083 = (f1083 >= `INH(p1030)) ? `INH(p1030) : f1083;
        f1084 = 4095;
        f1084 = (f1084 >= `INH(p1030)) ? `INH(p1030) : f1084;
        f1084 = (f1084 > p1031) ? p1031 : f1084;
        f1085 = 4095;
        f1085 = (f1085 > p1029) ? p1029 : f1085;
        f1085 = (f1085 >= `INH(p1031)) ? `INH(p1031) : f1085;
        f1086 = 4095;
        f1086 = (f1086 > p1019) ? p1019 : f1086;
        f1086 = (f1086 > p1026) ? p1026 : f1086;
        f1086 = (f1086 >= `INH(p1027)) ? `INH(p1027) : f1086;
        f1086 = (f1086 >= `INH(p1031)) ? `INH(p1031) : f1086;
        f1087 = 4095;
        f1087 = (f1087 > p1019) ? p1019 : f1087;
        f1087 = (f1087 >= `INH(p1026)) ? `INH(p1026) : f1087;
        f1087 = (f1087 >= `INH(p1031)) ? `INH(p1031) : f1087;
        f1088 = 4095;
        f1088 = (f1088 > p151) ? p151 : f1088;
        f1088 = (f1088 >= `INH(p1033)) ? `INH(p1033) : f1088;
        f1089 = 4095;
        f1089 = (f1089 > p1032) ? p1032 : f1089;
        f1089 = (f1089 >= `INH(p1034)) ? `INH(p1034) : f1089;
        f1090 = 4095;
        f1090 = (f1090 >= `INH(p151)) ? `INH(p151) : f1090;
        f1090 = (f1090 >= `INH(p1033)) ? `INH(p1033) : f1090;
        f1090 = (f1090 > p1034) ? p1034 : f1090;
        f1091 = 4095;
        f1091 = (f1091 >= `INH(p1032)) ? `INH(p1032) : f1091;
        f1091 = (f1091 >= `INH(p1034)) ? `INH(p1034) : f1091;
        f1091 = (f1091 > p1035) ? p1035 : f1091;
        f1092 = 4095;
        f1092 = (f1092 > p152) ? p152 : f1092;
        f1092 = (f1092 >= `INH(p1037)) ? `INH(p1037) : f1092;
        f1093 = 4095;
        f1093 = (f1093 > p1036) ? p1036 : f1093;
        f1093 = (f1093 >= `INH(p1038)) ? `INH(p1038) : f1093;
        f1094 = 4095;
        f1094 = (f1094 >= `INH(p152)) ? `INH(p152) : f1094;
        f1094 = (f1094 >= `INH(p1037)) ? `INH(p1037) : f1094;
        f1094 = (f1094 > p1038) ? p1038 : f1094;
        f1095 = 4095;
        f1095 = (f1095 >= `INH(p1036)) ? `INH(p1036) : f1095;
        f1095 = (f1095 >= `INH(p1038)) ? `INH(p1038) : f1095;
        f1095 = (f1095 > p1039) ? p1039 : f1095;
        f1096 = 4095;
        f1096 = (f1096 >= `INH(p141)) ? `INH(p141) : f1096;
        f1096 = (f1096 > p1033) ? p1033 : f1096;
        f1096 = (f1096 > p1037) ? p1037 : f1096;
        f1097 = 4095;
        f1097 = (f1097 > p1019) ? p1019 : f1097;
        f1097 = (f1097 >= `INH(p1035)) ? `INH(p1035) : f1097;
        f1097 = (f1097 >= `INH(p1039)) ? `INH(p1039) : f1097;
        f1098 = 4095;
        f1098 = (f1098 > p1020) ? p1020 : f1098;
        f1098 = (f1098 >= `INH(p1040)) ? `INH(p1040) : f1098;
        f1099 = 4095;
        f1099 = (f1099 > p153) ? p153 : f1099;
        f1099 = (f1099 >= `INH(p1021)) ? `INH(p1021) : f1099;
        f1100 = 4095;
        f1100 = (f1100 >= `INH(p153)) ? `INH(p153) : f1100;
        f1100 = (f1100 >= `INH(p1021)) ? `INH(p1021) : f1100;
        f1100 = (f1100 > p1040) ? p1040 : f1100;
        f1101 = 4095;
        f1101 = (f1101 > p142) ? p142 : f1101;
        f1101 = (f1101 >= `INH(p1020)) ? `INH(p1020) : f1101;
        f1101 = (f1101 >= `INH(p1040)) ? `INH(p1040) : f1101;
        f1102 = 4095;
        f1102 = (f1102 > p1042) ? p1042 : f1102;
        f1102 = (f1102 >= `INH(p1044)) ? `INH(p1044) : f1102;
        f1103 = 4095;
        f1103 = (f1103 >= `INH(p1041)) ? `INH(p1041) : f1103;
        f1103 = (f1103 >= `INH(p1042)) ? `INH(p1042) : f1103;
        f1103 = (f1103 >= `INH(p1044)) ? `INH(p1044) : f1103;
        f1103 = (f1103 > p1045) ? p1045 : f1103;
        f1104 = 4095;
        f1104 = (f1104 > p150) ? p150 : f1104;
        f1104 = (f1104 >= `INH(p1047)) ? `INH(p1047) : f1104;
        f1105 = 4095;
        f1105 = (f1105 > p1046) ? p1046 : f1105;
        f1105 = (f1105 >= `INH(p1048)) ? `INH(p1048) : f1105;
        f1106 = 4095;
        f1106 = (f1106 >= `INH(p150)) ? `INH(p150) : f1106;
        f1106 = (f1106 >= `INH(p1047)) ? `INH(p1047) : f1106;
        f1106 = (f1106 > p1048) ? p1048 : f1106;
        f1107 = 4095;
        f1107 = (f1107 >= `INH(p1046)) ? `INH(p1046) : f1107;
        f1107 = (f1107 >= `INH(p1048)) ? `INH(p1048) : f1107;
        f1107 = (f1107 > p1049) ? p1049 : f1107;
        f1108 = 4095;
        f1108 = (f1108 > p153) ? p153 : f1108;
        f1108 = (f1108 >= `INH(p1051)) ? `INH(p1051) : f1108;
        f1109 = 4095;
        f1109 = (f1109 > p1050) ? p1050 : f1109;
        f1109 = (f1109 >= `INH(p1052)) ? `INH(p1052) : f1109;
        f1110 = 4095;
        f1110 = (f1110 >= `INH(p153)) ? `INH(p153) : f1110;
        f1110 = (f1110 >= `INH(p1051)) ? `INH(p1051) : f1110;
        f1110 = (f1110 > p1052) ? p1052 : f1110;
        f1111 = 4095;
        f1111 = (f1111 >= `INH(p1050)) ? `INH(p1050) : f1111;
        f1111 = (f1111 >= `INH(p1052)) ? `INH(p1052) : f1111;
        f1111 = (f1111 > p1053) ? p1053 : f1111;
        f1112 = 4095;
        f1112 = (f1112 >= `INH(p142)) ? `INH(p142) : f1112;
        f1112 = (f1112 > p1047) ? p1047 : f1112;
        f1112 = (f1112 > p1051) ? p1051 : f1112;
        f1113 = 4095;
        f1113 = (f1113 > p1044) ? p1044 : f1113;
        f1113 = (f1113 >= `INH(p1049)) ? `INH(p1049) : f1113;
        f1113 = (f1113 >= `INH(p1053)) ? `INH(p1053) : f1113;
        f1114 = 4095;
        f1114 = (f1114 > p1043) ? p1043 : f1114;
        f1114 = (f1114 >= `INH(p1054)) ? `INH(p1054) : f1114;
        f1115 = 4095;
        f1115 = (f1115 > p154) ? p154 : f1115;
        f1115 = (f1115 >= `INH(p1045)) ? `INH(p1045) : f1115;
        f1116 = 4095;
        f1116 = (f1116 >= `INH(p154)) ? `INH(p154) : f1116;
        f1116 = (f1116 >= `INH(p1045)) ? `INH(p1045) : f1116;
        f1116 = (f1116 > p1054) ? p1054 : f1116;
        f1117 = 4095;
        f1117 = (f1117 > p143) ? p143 : f1117;
        f1117 = (f1117 >= `INH(p1043)) ? `INH(p1043) : f1117;
        f1117 = (f1117 >= `INH(p1054)) ? `INH(p1054) : f1117;
        if(f47>0)
                f2 = 0;
        if(f48>0)
                f49 = 0;
        if(f50>0)
                f51 = 0;
        if(f52>0)
                f53 = 0;
        if(f54>0)
                f56 = 0;
        if(f55>0)
                f56 = 0;
        if(f57>0)
                f58 = 0;
        if(f59>0)
                f60 = 0;
        if(f59>0)
                f61 = 0;
        if(f76>0)
                f3 = 0;
        if(f77>0)
                f78 = 0;
        if(f79>0)
                f80 = 0;
        if(f81>0)
                f82 = 0;
        if(f83>0)
                f85 = 0;
        if(f84>0)
                f85 = 0;
        if(f86>0)
                f87 = 0;
        if(f88>0)
                f89 = 0;
        if(f88>0)
                f90 = 0;
        if(f121>0)
                f5 = 0;
        if(f122>0)
                f123 = 0;
        if(f124>0)
                f125 = 0;
        if(f126>0)
                f127 = 0;
        if(f128>0)
                f130 = 0;
        if(f129>0)
                f130 = 0;
        if(f131>0)
                f132 = 0;
        if(f133>0)
                f134 = 0;
        if(f133>0)
                f135 = 0;
        if(f166>0)
                f7 = 0;
        if(f167>0)
                f168 = 0;
        if(f169>0)
                f170 = 0;
        if(f171>0)
                f172 = 0;
        if(f173>0)
                f175 = 0;
        if(f174>0)
                f175 = 0;
        if(f176>0)
                f177 = 0;
        if(f178>0)
                f179 = 0;
        if(f178>0)
                f180 = 0;
        if(f195>0)
                f8 = 0;
        if(f196>0)
                f197 = 0;
        if(f198>0)
                f199 = 0;
        if(f200>0)
                f201 = 0;
        if(f202>0)
                f204 = 0;
        if(f203>0)
                f204 = 0;
        if(f205>0)
                f206 = 0;
        if(f207>0)
                f208 = 0;
        if(f207>0)
                f209 = 0;
        if(f240>0)
                f10 = 0;
        if(f241>0)
                f242 = 0;
        if(f243>0)
                f244 = 0;
        if(f245>0)
                f246 = 0;
        if(f247>0)
                f249 = 0;
        if(f248>0)
                f249 = 0;
        if(f250>0)
                f251 = 0;
        if(f252>0)
                f253 = 0;
        if(f252>0)
                f254 = 0;
        if(f285>0)
                f12 = 0;
        if(f286>0)
                f287 = 0;
        if(f288>0)
                f289 = 0;
        if(f290>0)
                f291 = 0;
        if(f292>0)
                f294 = 0;
        if(f293>0)
                f294 = 0;
        if(f295>0)
                f296 = 0;
        if(f297>0)
                f298 = 0;
        if(f297>0)
                f299 = 0;
        if(f314>0)
                f13 = 0;
        if(f315>0)
                f316 = 0;
        if(f317>0)
                f318 = 0;
        if(f319>0)
                f320 = 0;
        if(f321>0)
                f323 = 0;
        if(f322>0)
                f323 = 0;
        if(f324>0)
                f325 = 0;
        if(f326>0)
                f327 = 0;
        if(f326>0)
                f328 = 0;
        if(f359>0)
                f15 = 0;
        if(f360>0)
                f361 = 0;
        if(f362>0)
                f363 = 0;
        if(f364>0)
                f365 = 0;
        if(f366>0)
                f368 = 0;
        if(f367>0)
                f368 = 0;
        if(f369>0)
                f370 = 0;
        if(f371>0)
                f372 = 0;
        if(f371>0)
                f373 = 0;
        if(f404>0)
                f17 = 0;
        if(f405>0)
                f406 = 0;
        if(f407>0)
                f408 = 0;
        if(f409>0)
                f410 = 0;
        if(f411>0)
                f413 = 0;
        if(f412>0)
                f413 = 0;
        if(f414>0)
                f415 = 0;
        if(f416>0)
                f417 = 0;
        if(f416>0)
                f418 = 0;
        if(f433>0)
                f18 = 0;
        if(f434>0)
                f435 = 0;
        if(f436>0)
                f437 = 0;
        if(f438>0)
                f439 = 0;
        if(f440>0)
                f442 = 0;
        if(f441>0)
                f442 = 0;
        if(f443>0)
                f444 = 0;
        if(f445>0)
                f446 = 0;
        if(f445>0)
                f447 = 0;
        if(f478>0)
                f20 = 0;
        if(f479>0)
                f480 = 0;
        if(f481>0)
                f482 = 0;
        if(f483>0)
                f484 = 0;
        if(f485>0)
                f487 = 0;
        if(f486>0)
                f487 = 0;
        if(f488>0)
                f489 = 0;
        if(f490>0)
                f491 = 0;
        if(f490>0)
                f492 = 0;
        if(f523>0)
                f22 = 0;
        if(f524>0)
                f525 = 0;
        if(f526>0)
                f527 = 0;
        if(f528>0)
                f529 = 0;
        if(f530>0)
                f532 = 0;
        if(f531>0)
                f532 = 0;
        if(f533>0)
                f534 = 0;
        if(f535>0)
                f536 = 0;
        if(f535>0)
                f537 = 0;
        if(f552>0)
                f23 = 0;
        if(f553>0)
                f554 = 0;
        if(f555>0)
                f556 = 0;
        if(f557>0)
                f558 = 0;
        if(f559>0)
                f561 = 0;
        if(f560>0)
                f561 = 0;
        if(f562>0)
                f563 = 0;
        if(f564>0)
                f565 = 0;
        if(f564>0)
                f566 = 0;
        if(f597>0)
                f25 = 0;
        if(f598>0)
                f599 = 0;
        if(f600>0)
                f601 = 0;
        if(f602>0)
                f603 = 0;
        if(f604>0)
                f606 = 0;
        if(f605>0)
                f606 = 0;
        if(f607>0)
                f608 = 0;
        if(f609>0)
                f610 = 0;
        if(f609>0)
                f611 = 0;
        if(f642>0)
                f27 = 0;
        if(f643>0)
                f644 = 0;
        if(f645>0)
                f646 = 0;
        if(f647>0)
                f648 = 0;
        if(f649>0)
                f651 = 0;
        if(f650>0)
                f651 = 0;
        if(f652>0)
                f653 = 0;
        if(f654>0)
                f655 = 0;
        if(f654>0)
                f656 = 0;
        if(f671>0)
                f28 = 0;
        if(f672>0)
                f673 = 0;
        if(f674>0)
                f675 = 0;
        if(f676>0)
                f677 = 0;
        if(f678>0)
                f680 = 0;
        if(f679>0)
                f680 = 0;
        if(f681>0)
                f682 = 0;
        if(f683>0)
                f684 = 0;
        if(f683>0)
                f685 = 0;
        if(f716>0)
                f30 = 0;
        if(f717>0)
                f718 = 0;
        if(f719>0)
                f720 = 0;
        if(f721>0)
                f722 = 0;
        if(f723>0)
                f725 = 0;
        if(f724>0)
                f725 = 0;
        if(f726>0)
                f727 = 0;
        if(f728>0)
                f729 = 0;
        if(f728>0)
                f730 = 0;
        if(f761>0)
                f32 = 0;
        if(f762>0)
                f763 = 0;
        if(f764>0)
                f765 = 0;
        if(f766>0)
                f767 = 0;
        if(f768>0)
                f770 = 0;
        if(f769>0)
                f770 = 0;
        if(f771>0)
                f772 = 0;
        if(f773>0)
                f774 = 0;
        if(f773>0)
                f775 = 0;
        if(f790>0)
                f33 = 0;
        if(f791>0)
                f792 = 0;
        if(f793>0)
                f794 = 0;
        if(f795>0)
                f796 = 0;
        if(f797>0)
                f799 = 0;
        if(f798>0)
                f799 = 0;
        if(f800>0)
                f801 = 0;
        if(f802>0)
                f803 = 0;
        if(f802>0)
                f804 = 0;
        if(f835>0)
                f35 = 0;
        if(f836>0)
                f837 = 0;
        if(f838>0)
                f839 = 0;
        if(f840>0)
                f841 = 0;
        if(f842>0)
                f844 = 0;
        if(f843>0)
                f844 = 0;
        if(f845>0)
                f846 = 0;
        if(f847>0)
                f848 = 0;
        if(f847>0)
                f849 = 0;
        if(f880>0)
                f37 = 0;
        if(f881>0)
                f882 = 0;
        if(f883>0)
                f884 = 0;
        if(f885>0)
                f886 = 0;
        if(f887>0)
                f889 = 0;
        if(f888>0)
                f889 = 0;
        if(f890>0)
                f891 = 0;
        if(f892>0)
                f893 = 0;
        if(f892>0)
                f894 = 0;
        if(f909>0)
                f38 = 0;
        if(f910>0)
                f911 = 0;
        if(f912>0)
                f913 = 0;
        if(f914>0)
                f915 = 0;
        if(f916>0)
                f918 = 0;
        if(f917>0)
                f918 = 0;
        if(f919>0)
                f920 = 0;
        if(f921>0)
                f922 = 0;
        if(f921>0)
                f923 = 0;
        if(f954>0)
                f40 = 0;
        if(f955>0)
                f956 = 0;
        if(f957>0)
                f958 = 0;
        if(f959>0)
                f960 = 0;
        if(f961>0)
                f963 = 0;
        if(f962>0)
                f963 = 0;
        if(f964>0)
                f965 = 0;
        if(f966>0)
                f967 = 0;
        if(f966>0)
                f968 = 0;
        if(f999>0)
                f42 = 0;
        if(f1000>0)
                f1001 = 0;
        if(f1002>0)
                f1003 = 0;
        if(f1004>0)
                f1005 = 0;
        if(f1006>0)
                f1008 = 0;
        if(f1007>0)
                f1008 = 0;
        if(f1009>0)
                f1010 = 0;
        if(f1011>0)
                f1012 = 0;
        if(f1011>0)
                f1013 = 0;
        if(f1028>0)
                f43 = 0;
        if(f1029>0)
                f1030 = 0;
        if(f1031>0)
                f1032 = 0;
        if(f1033>0)
                f1034 = 0;
        if(f1035>0)
                f1037 = 0;
        if(f1036>0)
                f1037 = 0;
        if(f1038>0)
                f1039 = 0;
        if(f1040>0)
                f1041 = 0;
        if(f1040>0)
                f1042 = 0;
        if(f1073>0)
                f45 = 0;
        if(f1074>0)
                f1075 = 0;
        if(f1076>0)
                f1077 = 0;
        if(f1078>0)
                f1079 = 0;
        if(f1080>0)
                f1082 = 0;
        if(f1081>0)
                f1082 = 0;
        if(f1083>0)
                f1084 = 0;
        if(f1085>0)
                f1086 = 0;
        if(f1085>0)
                f1087 = 0;
        tf = (f0>0)?1:(f1>0)?2:(f2>0)?3:(f3>0)?4:(f4>0)?5:(f5>0)?6:(f6>0)?7:(f7>0)?8:(f8>0)?9:(f9>0)?10:(f10>0)?11:(f11>0)?12:(f12>0)?13:(f13>0)?14:(f14>0)?15:(f15>0)?16:(f16>0)?17:(f17>0)?18:(f18>0)?19:(f19>0)?20:(f20>0)?21:(f21>0)?22:(f22>0)?23:(f23>0)?24:(f24>0)?25:(f25>0)?26:(f26>0)?27:(f27>0)?28:(f28>0)?29:(f29>0)?30:(f30>0)?31:(f31>0)?32:(f32>0)?33:(f33>0)?34:(f34>0)?35:(f35>0)?36:(f36>0)?37:(f37>0)?38:(f38>0)?39:(f39>0)?40:(f40>0)?41:(f41>0)?42:(f42>0)?43:(f43>0)?44:(f44>0)?45:(f45>0)?46:(f46>0)?47:(f47>0)?48:(f48>0)?49:(f49>0)?50:(f50>0)?51:(f51>0)?52:(f52>0)?53:(f53>0)?54:(f54>0)?55:(f55>0)?56:(f56>0)?57:(f57>0)?58:(f58>0)?59:(f59>0)?60:(f60>0)?61:(f61>0)?62:(f62>0)?63:(f63>0)?64:(f64>0)?65:(f65>0)?66:(f66>0)?67:(f67>0)?68:(f68>0)?69:(f69>0)?70:(f70>0)?71:(f71>0)?72:(f72>0)?73:(f73>0)?74:(f74>0)?75:(f75>0)?76:(f76>0)?77:(f77>0)?78:(f78>0)?79:(f79>0)?80:(f80>0)?81:(f81>0)?82:(f82>0)?83:(f83>0)?84:(f84>0)?85:(f85>0)?86:(f86>0)?87:(f87>0)?88:(f88>0)?89:(f89>0)?90:(f90>0)?91:(f91>0)?92:(f92>0)?93:(f93>0)?94:(f94>0)?95:(f95>0)?96:(f96>0)?97:(f97>0)?98:(f98>0)?99:(f99>0)?100:(f100>0)?101:(f101>0)?102:(f102>0)?103:(f103>0)?104:(f104>0)?105:(f105>0)?106:(f106>0)?107:(f107>0)?108:(f108>0)?109:(f109>0)?110:(f110>0)?111:(f111>0)?112:(f112>0)?113:(f113>0)?114:(f114>0)?115:(f115>0)?116:(f116>0)?117:(f117>0)?118:(f118>0)?119:(f119>0)?120:(f120>0)?121:(f121>0)?122:(f122>0)?123:(f123>0)?124:(f124>0)?125:(f125>0)?126:(f126>0)?127:(f127>0)?128:(f128>0)?129:(f129>0)?130:(f130>0)?131:(f131>0)?132:(f132>0)?133:(f133>0)?134:(f134>0)?135:(f135>0)?136:(f136>0)?137:(f137>0)?138:(f138>0)?139:(f139>0)?140:(f140>0)?141:(f141>0)?142:(f142>0)?143:(f143>0)?144:(f144>0)?145:(f145>0)?146:(f146>0)?147:(f147>0)?148:(f148>0)?149:(f149>0)?150:(f150>0)?151:(f151>0)?152:(f152>0)?153:(f153>0)?154:(f154>0)?155:(f155>0)?156:(f156>0)?157:(f157>0)?158:(f158>0)?159:(f159>0)?160:(f160>0)?161:(f161>0)?162:(f162>0)?163:(f163>0)?164:(f164>0)?165:(f165>0)?166:(f166>0)?167:(f167>0)?168:(f168>0)?169:(f169>0)?170:(f170>0)?171:(f171>0)?172:(f172>0)?173:(f173>0)?174:(f174>0)?175:(f175>0)?176:(f176>0)?177:(f177>0)?178:(f178>0)?179:(f179>0)?180:(f180>0)?181:(f181>0)?182:(f182>0)?183:(f183>0)?184:(f184>0)?185:(f185>0)?186:(f186>0)?187:(f187>0)?188:(f188>0)?189:(f189>0)?190:(f190>0)?191:(f191>0)?192:(f192>0)?193:(f193>0)?194:(f194>0)?195:(f195>0)?196:(f196>0)?197:(f197>0)?198:(f198>0)?199:(f199>0)?200:(f200>0)?201:(f201>0)?202:(f202>0)?203:(f203>0)?204:(f204>0)?205:(f205>0)?206:(f206>0)?207:(f207>0)?208:(f208>0)?209:(f209>0)?210:(f210>0)?211:(f211>0)?212:(f212>0)?213:(f213>0)?214:(f214>0)?215:(f215>0)?216:(f216>0)?217:(f217>0)?218:(f218>0)?219:(f219>0)?220:(f220>0)?221:(f221>0)?222:(f222>0)?223:(f223>0)?224:(f224>0)?225:(f225>0)?226:(f226>0)?227:(f227>0)?228:(f228>0)?229:(f229>0)?230:(f230>0)?231:(f231>0)?232:(f232>0)?233:(f233>0)?234:(f234>0)?235:(f235>0)?236:(f236>0)?237:(f237>0)?238:(f238>0)?239:(f239>0)?240:(f240>0)?241:(f241>0)?242:(f242>0)?243:(f243>0)?244:(f244>0)?245:(f245>0)?246:(f246>0)?247:(f247>0)?248:(f248>0)?249:(f249>0)?250:(f250>0)?251:(f251>0)?252:(f252>0)?253:(f253>0)?254:(f254>0)?255:(f255>0)?256:(f256>0)?257:(f257>0)?258:(f258>0)?259:(f259>0)?260:(f260>0)?261:(f261>0)?262:(f262>0)?263:(f263>0)?264:(f264>0)?265:(f265>0)?266:(f266>0)?267:(f267>0)?268:(f268>0)?269:(f269>0)?270:(f270>0)?271:(f271>0)?272:(f272>0)?273:(f273>0)?274:(f274>0)?275:(f275>0)?276:(f276>0)?277:(f277>0)?278:(f278>0)?279:(f279>0)?280:(f280>0)?281:(f281>0)?282:(f282>0)?283:(f283>0)?284:(f284>0)?285:(f285>0)?286:(f286>0)?287:(f287>0)?288:(f288>0)?289:(f289>0)?290:(f290>0)?291:(f291>0)?292:(f292>0)?293:(f293>0)?294:(f294>0)?295:(f295>0)?296:(f296>0)?297:(f297>0)?298:(f298>0)?299:(f299>0)?300:(f300>0)?301:(f301>0)?302:(f302>0)?303:(f303>0)?304:(f304>0)?305:(f305>0)?306:(f306>0)?307:(f307>0)?308:(f308>0)?309:(f309>0)?310:(f310>0)?311:(f311>0)?312:(f312>0)?313:(f313>0)?314:(f314>0)?315:(f315>0)?316:(f316>0)?317:(f317>0)?318:(f318>0)?319:(f319>0)?320:(f320>0)?321:(f321>0)?322:(f322>0)?323:(f323>0)?324:(f324>0)?325:(f325>0)?326:(f326>0)?327:(f327>0)?328:(f328>0)?329:(f329>0)?330:(f330>0)?331:(f331>0)?332:(f332>0)?333:(f333>0)?334:(f334>0)?335:(f335>0)?336:(f336>0)?337:(f337>0)?338:(f338>0)?339:(f339>0)?340:(f340>0)?341:(f341>0)?342:(f342>0)?343:(f343>0)?344:(f344>0)?345:(f345>0)?346:(f346>0)?347:(f347>0)?348:(f348>0)?349:(f349>0)?350:(f350>0)?351:(f351>0)?352:(f352>0)?353:(f353>0)?354:(f354>0)?355:(f355>0)?356:(f356>0)?357:(f357>0)?358:(f358>0)?359:(f359>0)?360:(f360>0)?361:(f361>0)?362:(f362>0)?363:(f363>0)?364:(f364>0)?365:(f365>0)?366:(f366>0)?367:(f367>0)?368:(f368>0)?369:(f369>0)?370:(f370>0)?371:(f371>0)?372:(f372>0)?373:(f373>0)?374:(f374>0)?375:(f375>0)?376:(f376>0)?377:(f377>0)?378:(f378>0)?379:(f379>0)?380:(f380>0)?381:(f381>0)?382:(f382>0)?383:(f383>0)?384:(f384>0)?385:(f385>0)?386:(f386>0)?387:(f387>0)?388:(f388>0)?389:(f389>0)?390:(f390>0)?391:(f391>0)?392:(f392>0)?393:(f393>0)?394:(f394>0)?395:(f395>0)?396:(f396>0)?397:(f397>0)?398:(f398>0)?399:(f399>0)?400:(f400>0)?401:(f401>0)?402:(f402>0)?403:(f403>0)?404:(f404>0)?405:(f405>0)?406:(f406>0)?407:(f407>0)?408:(f408>0)?409:(f409>0)?410:(f410>0)?411:(f411>0)?412:(f412>0)?413:(f413>0)?414:(f414>0)?415:(f415>0)?416:(f416>0)?417:(f417>0)?418:(f418>0)?419:(f419>0)?420:(f420>0)?421:(f421>0)?422:(f422>0)?423:(f423>0)?424:(f424>0)?425:(f425>0)?426:(f426>0)?427:(f427>0)?428:(f428>0)?429:(f429>0)?430:(f430>0)?431:(f431>0)?432:(f432>0)?433:(f433>0)?434:(f434>0)?435:(f435>0)?436:(f436>0)?437:(f437>0)?438:(f438>0)?439:(f439>0)?440:(f440>0)?441:(f441>0)?442:(f442>0)?443:(f443>0)?444:(f444>0)?445:(f445>0)?446:(f446>0)?447:(f447>0)?448:(f448>0)?449:(f449>0)?450:(f450>0)?451:(f451>0)?452:(f452>0)?453:(f453>0)?454:(f454>0)?455:(f455>0)?456:(f456>0)?457:(f457>0)?458:(f458>0)?459:(f459>0)?460:(f460>0)?461:(f461>0)?462:(f462>0)?463:(f463>0)?464:(f464>0)?465:(f465>0)?466:(f466>0)?467:(f467>0)?468:(f468>0)?469:(f469>0)?470:(f470>0)?471:(f471>0)?472:(f472>0)?473:(f473>0)?474:(f474>0)?475:(f475>0)?476:(f476>0)?477:(f477>0)?478:(f478>0)?479:(f479>0)?480:(f480>0)?481:(f481>0)?482:(f482>0)?483:(f483>0)?484:(f484>0)?485:(f485>0)?486:(f486>0)?487:(f487>0)?488:(f488>0)?489:(f489>0)?490:(f490>0)?491:(f491>0)?492:(f492>0)?493:(f493>0)?494:(f494>0)?495:(f495>0)?496:(f496>0)?497:(f497>0)?498:(f498>0)?499:(f499>0)?500:(f500>0)?501:(f501>0)?502:(f502>0)?503:(f503>0)?504:(f504>0)?505:(f505>0)?506:(f506>0)?507:(f507>0)?508:(f508>0)?509:(f509>0)?510:(f510>0)?511:(f511>0)?512:(f512>0)?513:(f513>0)?514:(f514>0)?515:(f515>0)?516:(f516>0)?517:(f517>0)?518:(f518>0)?519:(f519>0)?520:(f520>0)?521:(f521>0)?522:(f522>0)?523:(f523>0)?524:(f524>0)?525:(f525>0)?526:(f526>0)?527:(f527>0)?528:(f528>0)?529:(f529>0)?530:(f530>0)?531:(f531>0)?532:(f532>0)?533:(f533>0)?534:(f534>0)?535:(f535>0)?536:(f536>0)?537:(f537>0)?538:(f538>0)?539:(f539>0)?540:(f540>0)?541:(f541>0)?542:(f542>0)?543:(f543>0)?544:(f544>0)?545:(f545>0)?546:(f546>0)?547:(f547>0)?548:(f548>0)?549:(f549>0)?550:(f550>0)?551:(f551>0)?552:(f552>0)?553:(f553>0)?554:(f554>0)?555:(f555>0)?556:(f556>0)?557:(f557>0)?558:(f558>0)?559:(f559>0)?560:(f560>0)?561:(f561>0)?562:(f562>0)?563:(f563>0)?564:(f564>0)?565:(f565>0)?566:(f566>0)?567:(f567>0)?568:(f568>0)?569:(f569>0)?570:(f570>0)?571:(f571>0)?572:(f572>0)?573:(f573>0)?574:(f574>0)?575:(f575>0)?576:(f576>0)?577:(f577>0)?578:(f578>0)?579:(f579>0)?580:(f580>0)?581:(f581>0)?582:(f582>0)?583:(f583>0)?584:(f584>0)?585:(f585>0)?586:(f586>0)?587:(f587>0)?588:(f588>0)?589:(f589>0)?590:(f590>0)?591:(f591>0)?592:(f592>0)?593:(f593>0)?594:(f594>0)?595:(f595>0)?596:(f596>0)?597:(f597>0)?598:(f598>0)?599:(f599>0)?600:(f600>0)?601:(f601>0)?602:(f602>0)?603:(f603>0)?604:(f604>0)?605:(f605>0)?606:(f606>0)?607:(f607>0)?608:(f608>0)?609:(f609>0)?610:(f610>0)?611:(f611>0)?612:(f612>0)?613:(f613>0)?614:(f614>0)?615:(f615>0)?616:(f616>0)?617:(f617>0)?618:(f618>0)?619:(f619>0)?620:(f620>0)?621:(f621>0)?622:(f622>0)?623:(f623>0)?624:(f624>0)?625:(f625>0)?626:(f626>0)?627:(f627>0)?628:(f628>0)?629:(f629>0)?630:(f630>0)?631:(f631>0)?632:(f632>0)?633:(f633>0)?634:(f634>0)?635:(f635>0)?636:(f636>0)?637:(f637>0)?638:(f638>0)?639:(f639>0)?640:(f640>0)?641:(f641>0)?642:(f642>0)?643:(f643>0)?644:(f644>0)?645:(f645>0)?646:(f646>0)?647:(f647>0)?648:(f648>0)?649:(f649>0)?650:(f650>0)?651:(f651>0)?652:(f652>0)?653:(f653>0)?654:(f654>0)?655:(f655>0)?656:(f656>0)?657:(f657>0)?658:(f658>0)?659:(f659>0)?660:(f660>0)?661:(f661>0)?662:(f662>0)?663:(f663>0)?664:(f664>0)?665:(f665>0)?666:(f666>0)?667:(f667>0)?668:(f668>0)?669:(f669>0)?670:(f670>0)?671:(f671>0)?672:(f672>0)?673:(f673>0)?674:(f674>0)?675:(f675>0)?676:(f676>0)?677:(f677>0)?678:(f678>0)?679:(f679>0)?680:(f680>0)?681:(f681>0)?682:(f682>0)?683:(f683>0)?684:(f684>0)?685:(f685>0)?686:(f686>0)?687:(f687>0)?688:(f688>0)?689:(f689>0)?690:(f690>0)?691:(f691>0)?692:(f692>0)?693:(f693>0)?694:(f694>0)?695:(f695>0)?696:(f696>0)?697:(f697>0)?698:(f698>0)?699:(f699>0)?700:(f700>0)?701:(f701>0)?702:(f702>0)?703:(f703>0)?704:(f704>0)?705:(f705>0)?706:(f706>0)?707:(f707>0)?708:(f708>0)?709:(f709>0)?710:(f710>0)?711:(f711>0)?712:(f712>0)?713:(f713>0)?714:(f714>0)?715:(f715>0)?716:(f716>0)?717:(f717>0)?718:(f718>0)?719:(f719>0)?720:(f720>0)?721:(f721>0)?722:(f722>0)?723:(f723>0)?724:(f724>0)?725:(f725>0)?726:(f726>0)?727:(f727>0)?728:(f728>0)?729:(f729>0)?730:(f730>0)?731:(f731>0)?732:(f732>0)?733:(f733>0)?734:(f734>0)?735:(f735>0)?736:(f736>0)?737:(f737>0)?738:(f738>0)?739:(f739>0)?740:(f740>0)?741:(f741>0)?742:(f742>0)?743:(f743>0)?744:(f744>0)?745:(f745>0)?746:(f746>0)?747:(f747>0)?748:(f748>0)?749:(f749>0)?750:(f750>0)?751:(f751>0)?752:(f752>0)?753:(f753>0)?754:(f754>0)?755:(f755>0)?756:(f756>0)?757:(f757>0)?758:(f758>0)?759:(f759>0)?760:(f760>0)?761:(f761>0)?762:(f762>0)?763:(f763>0)?764:(f764>0)?765:(f765>0)?766:(f766>0)?767:(f767>0)?768:(f768>0)?769:(f769>0)?770:(f770>0)?771:(f771>0)?772:(f772>0)?773:(f773>0)?774:(f774>0)?775:(f775>0)?776:(f776>0)?777:(f777>0)?778:(f778>0)?779:(f779>0)?780:(f780>0)?781:(f781>0)?782:(f782>0)?783:(f783>0)?784:(f784>0)?785:(f785>0)?786:(f786>0)?787:(f787>0)?788:(f788>0)?789:(f789>0)?790:(f790>0)?791:(f791>0)?792:(f792>0)?793:(f793>0)?794:(f794>0)?795:(f795>0)?796:(f796>0)?797:(f797>0)?798:(f798>0)?799:(f799>0)?800:(f800>0)?801:(f801>0)?802:(f802>0)?803:(f803>0)?804:(f804>0)?805:(f805>0)?806:(f806>0)?807:(f807>0)?808:(f808>0)?809:(f809>0)?810:(f810>0)?811:(f811>0)?812:(f812>0)?813:(f813>0)?814:(f814>0)?815:(f815>0)?816:(f816>0)?817:(f817>0)?818:(f818>0)?819:(f819>0)?820:(f820>0)?821:(f821>0)?822:(f822>0)?823:(f823>0)?824:(f824>0)?825:(f825>0)?826:(f826>0)?827:(f827>0)?828:(f828>0)?829:(f829>0)?830:(f830>0)?831:(f831>0)?832:(f832>0)?833:(f833>0)?834:(f834>0)?835:(f835>0)?836:(f836>0)?837:(f837>0)?838:(f838>0)?839:(f839>0)?840:(f840>0)?841:(f841>0)?842:(f842>0)?843:(f843>0)?844:(f844>0)?845:(f845>0)?846:(f846>0)?847:(f847>0)?848:(f848>0)?849:(f849>0)?850:(f850>0)?851:(f851>0)?852:(f852>0)?853:(f853>0)?854:(f854>0)?855:(f855>0)?856:(f856>0)?857:(f857>0)?858:(f858>0)?859:(f859>0)?860:(f860>0)?861:(f861>0)?862:(f862>0)?863:(f863>0)?864:(f864>0)?865:(f865>0)?866:(f866>0)?867:(f867>0)?868:(f868>0)?869:(f869>0)?870:(f870>0)?871:(f871>0)?872:(f872>0)?873:(f873>0)?874:(f874>0)?875:(f875>0)?876:(f876>0)?877:(f877>0)?878:(f878>0)?879:(f879>0)?880:(f880>0)?881:(f881>0)?882:(f882>0)?883:(f883>0)?884:(f884>0)?885:(f885>0)?886:(f886>0)?887:(f887>0)?888:(f888>0)?889:(f889>0)?890:(f890>0)?891:(f891>0)?892:(f892>0)?893:(f893>0)?894:(f894>0)?895:(f895>0)?896:(f896>0)?897:(f897>0)?898:(f898>0)?899:(f899>0)?900:(f900>0)?901:(f901>0)?902:(f902>0)?903:(f903>0)?904:(f904>0)?905:(f905>0)?906:(f906>0)?907:(f907>0)?908:(f908>0)?909:(f909>0)?910:(f910>0)?911:(f911>0)?912:(f912>0)?913:(f913>0)?914:(f914>0)?915:(f915>0)?916:(f916>0)?917:(f917>0)?918:(f918>0)?919:(f919>0)?920:(f920>0)?921:(f921>0)?922:(f922>0)?923:(f923>0)?924:(f924>0)?925:(f925>0)?926:(f926>0)?927:(f927>0)?928:(f928>0)?929:(f929>0)?930:(f930>0)?931:(f931>0)?932:(f932>0)?933:(f933>0)?934:(f934>0)?935:(f935>0)?936:(f936>0)?937:(f937>0)?938:(f938>0)?939:(f939>0)?940:(f940>0)?941:(f941>0)?942:(f942>0)?943:(f943>0)?944:(f944>0)?945:(f945>0)?946:(f946>0)?947:(f947>0)?948:(f948>0)?949:(f949>0)?950:(f950>0)?951:(f951>0)?952:(f952>0)?953:(f953>0)?954:(f954>0)?955:(f955>0)?956:(f956>0)?957:(f957>0)?958:(f958>0)?959:(f959>0)?960:(f960>0)?961:(f961>0)?962:(f962>0)?963:(f963>0)?964:(f964>0)?965:(f965>0)?966:(f966>0)?967:(f967>0)?968:(f968>0)?969:(f969>0)?970:(f970>0)?971:(f971>0)?972:(f972>0)?973:(f973>0)?974:(f974>0)?975:(f975>0)?976:(f976>0)?977:(f977>0)?978:(f978>0)?979:(f979>0)?980:(f980>0)?981:(f981>0)?982:(f982>0)?983:(f983>0)?984:(f984>0)?985:(f985>0)?986:(f986>0)?987:(f987>0)?988:(f988>0)?989:(f989>0)?990:(f990>0)?991:(f991>0)?992:(f992>0)?993:(f993>0)?994:(f994>0)?995:(f995>0)?996:(f996>0)?997:(f997>0)?998:(f998>0)?999:(f999>0)?1000:(f1000>0)?1001:(f1001>0)?1002:(f1002>0)?1003:(f1003>0)?1004:(f1004>0)?1005:(f1005>0)?1006:(f1006>0)?1007:(f1007>0)?1008:(f1008>0)?1009:(f1009>0)?1010:(f1010>0)?1011:(f1011>0)?1012:(f1012>0)?1013:(f1013>0)?1014:(f1014>0)?1015:(f1015>0)?1016:(f1016>0)?1017:(f1017>0)?1018:(f1018>0)?1019:(f1019>0)?1020:(f1020>0)?1021:(f1021>0)?1022:(f1022>0)?1023:(f1023>0)?1024:(f1024>0)?1025:(f1025>0)?1026:(f1026>0)?1027:(f1027>0)?1028:(f1028>0)?1029:(f1029>0)?1030:(f1030>0)?1031:(f1031>0)?1032:(f1032>0)?1033:(f1033>0)?1034:(f1034>0)?1035:(f1035>0)?1036:(f1036>0)?1037:(f1037>0)?1038:(f1038>0)?1039:(f1039>0)?1040:(f1040>0)?1041:(f1041>0)?1042:(f1042>0)?1043:(f1043>0)?1044:(f1044>0)?1045:(f1045>0)?1046:(f1046>0)?1047:(f1047>0)?1048:(f1048>0)?1049:(f1049>0)?1050:(f1050>0)?1051:(f1051>0)?1052:(f1052>0)?1053:(f1053>0)?1054:(f1054>0)?1055:(f1055>0)?1056:(f1056>0)?1057:(f1057>0)?1058:(f1058>0)?1059:(f1059>0)?1060:(f1060>0)?1061:(f1061>0)?1062:(f1062>0)?1063:(f1063>0)?1064:(f1064>0)?1065:(f1065>0)?1066:(f1066>0)?1067:(f1067>0)?1068:(f1068>0)?1069:(f1069>0)?1070:(f1070>0)?1071:(f1071>0)?1072:(f1072>0)?1073:(f1073>0)?1074:(f1074>0)?1075:(f1075>0)?1076:(f1076>0)?1077:(f1077>0)?1078:(f1078>0)?1079:(f1079>0)?1080:(f1080>0)?1081:(f1081>0)?1082:(f1082>0)?1083:(f1083>0)?1084:(f1084>0)?1085:(f1085>0)?1086:(f1086>0)?1087:(f1087>0)?1088:(f1088>0)?1089:(f1089>0)?1090:(f1090>0)?1091:(f1091>0)?1092:(f1092>0)?1093:(f1093>0)?1094:(f1094>0)?1095:(f1095>0)?1096:(f1096>0)?1097:(f1097>0)?1098:(f1098>0)?1099:(f1099>0)?1100:(f1100>0)?1101:(f1101>0)?1102:(f1102>0)?1103:(f1103>0)?1104:(f1104>0)?1105:(f1105>0)?1106:(f1106>0)?1107:(f1107>0)?1108:(f1108>0)?1109:(f1109>0)?1110:(f1110>0)?1111:(f1111>0)?1112:(f1112>0)?1113:(f1113>0)?1114:(f1114>0)?1115:(f1115>0)?1116:(f1116>0)?1117:(f1117>0)?1118:0; 
       case(tf)
                1: begin
                        tc = f0;
                        p2 = p2 - tc;
                        p19 = p19 - tc;
                        p36 = p36 - tc;
                        p53 = p53 - tc;
                        p70 = p70 - tc;
                        p87 = p87 - tc;
                        p104 = p104 - tc;
                        p121 = p121 - tc;
                        p138 = p138 - tc;
                        p0 = p0 + tc;
                end
                2: begin
                        tc = f1;
                        p1 = p1 - tc;
                        p7 = p7 + tc;
                        p24 = p24 + tc;
                        p41 = p41 + tc;
                        p58 = p58 + tc;
                        p75 = p75 + tc;
                        p92 = p92 + tc;
                        p109 = p109 + tc;
                        p126 = p126 + tc;
                        p143 = p143 + tc;
                end
                3: begin
                        tc = f2;
                        p160 = p160 - tc;
                        p157 = p157 + tc;
                end
                4: begin
                        tc = f3;
                        p184 = p184 - tc;
                        p181 = p181 + tc;
                end
                5: begin
                        tc = f4;
                        p203 = p203 - tc;
                        p205 = p205 + tc;
                end
                6: begin
                        tc = f5;
                        p222 = p222 - tc;
                        p219 = p219 + tc;
                end
                7: begin
                        tc = f6;
                        p241 = p241 - tc;
                        p243 = p243 + tc;
                end
                8: begin
                        tc = f7;
                        p260 = p260 - tc;
                        p257 = p257 + tc;
                end
                9: begin
                        tc = f8;
                        p284 = p284 - tc;
                        p281 = p281 + tc;
                end
                10: begin
                        tc = f9;
                        p303 = p303 - tc;
                        p305 = p305 + tc;
                end
                11: begin
                        tc = f10;
                        p322 = p322 - tc;
                        p319 = p319 + tc;
                end
                12: begin
                        tc = f11;
                        p341 = p341 - tc;
                        p343 = p343 + tc;
                end
                13: begin
                        tc = f12;
                        p360 = p360 - tc;
                        p357 = p357 + tc;
                end
                14: begin
                        tc = f13;
                        p384 = p384 - tc;
                        p381 = p381 + tc;
                end
                15: begin
                        tc = f14;
                        p403 = p403 - tc;
                        p405 = p405 + tc;
                end
                16: begin
                        tc = f15;
                        p422 = p422 - tc;
                        p419 = p419 + tc;
                end
                17: begin
                        tc = f16;
                        p441 = p441 - tc;
                        p443 = p443 + tc;
                end
                18: begin
                        tc = f17;
                        p460 = p460 - tc;
                        p457 = p457 + tc;
                end
                19: begin
                        tc = f18;
                        p484 = p484 - tc;
                        p481 = p481 + tc;
                end
                20: begin
                        tc = f19;
                        p503 = p503 - tc;
                        p505 = p505 + tc;
                end
                21: begin
                        tc = f20;
                        p522 = p522 - tc;
                        p519 = p519 + tc;
                end
                22: begin
                        tc = f21;
                        p541 = p541 - tc;
                        p543 = p543 + tc;
                end
                23: begin
                        tc = f22;
                        p560 = p560 - tc;
                        p557 = p557 + tc;
                end
                24: begin
                        tc = f23;
                        p584 = p584 - tc;
                        p581 = p581 + tc;
                end
                25: begin
                        tc = f24;
                        p603 = p603 - tc;
                        p605 = p605 + tc;
                end
                26: begin
                        tc = f25;
                        p622 = p622 - tc;
                        p619 = p619 + tc;
                end
                27: begin
                        tc = f26;
                        p641 = p641 - tc;
                        p643 = p643 + tc;
                end
                28: begin
                        tc = f27;
                        p660 = p660 - tc;
                        p657 = p657 + tc;
                end
                29: begin
                        tc = f28;
                        p684 = p684 - tc;
                        p681 = p681 + tc;
                end
                30: begin
                        tc = f29;
                        p703 = p703 - tc;
                        p705 = p705 + tc;
                end
                31: begin
                        tc = f30;
                        p722 = p722 - tc;
                        p719 = p719 + tc;
                end
                32: begin
                        tc = f31;
                        p741 = p741 - tc;
                        p743 = p743 + tc;
                end
                33: begin
                        tc = f32;
                        p760 = p760 - tc;
                        p757 = p757 + tc;
                end
                34: begin
                        tc = f33;
                        p784 = p784 - tc;
                        p781 = p781 + tc;
                end
                35: begin
                        tc = f34;
                        p803 = p803 - tc;
                        p805 = p805 + tc;
                end
                36: begin
                        tc = f35;
                        p822 = p822 - tc;
                        p819 = p819 + tc;
                end
                37: begin
                        tc = f36;
                        p841 = p841 - tc;
                        p843 = p843 + tc;
                end
                38: begin
                        tc = f37;
                        p860 = p860 - tc;
                        p857 = p857 + tc;
                end
                39: begin
                        tc = f38;
                        p884 = p884 - tc;
                        p881 = p881 + tc;
                end
                40: begin
                        tc = f39;
                        p903 = p903 - tc;
                        p905 = p905 + tc;
                end
                41: begin
                        tc = f40;
                        p922 = p922 - tc;
                        p919 = p919 + tc;
                end
                42: begin
                        tc = f41;
                        p941 = p941 - tc;
                        p943 = p943 + tc;
                end
                43: begin
                        tc = f42;
                        p960 = p960 - tc;
                        p957 = p957 + tc;
                end
                44: begin
                        tc = f43;
                        p984 = p984 - tc;
                        p981 = p981 + tc;
                end
                45: begin
                        tc = f44;
                        p1003 = p1003 - tc;
                        p1005 = p1005 + tc;
                end
                46: begin
                        tc = f45;
                        p1022 = p1022 - tc;
                        p1019 = p1019 + tc;
                end
                47: begin
                        tc = f46;
                        p1041 = p1041 - tc;
                        p1043 = p1043 + tc;
                end
                48: begin
                        tc = f47;
                        p161 = p161 - tc;
                        p157 = p157 + tc;
                end
                49: begin
                        tc = f48;
                        p155 = p155 - tc;
                end
                50: begin
                        tc = f49;
                        p159 = p159 - tc;
                        p161 = p161 + tc;
                end
                51: begin
                        tc = f50;
                        p156 = p156 - tc*2;
                        p162 = p162 + tc;
                end
                52: begin
                        tc = f51;
                        p163 = p163 - tc;
                        p160 = p160 + tc;
                end
                53: begin
                        tc = f52;
                        p156 = p156 - tc;
                        p165 = p165 - tc;
                        p164 = p164 + tc;
                end
                54: begin
                        tc = f53;
                        p166 = p166 - tc;
                        p163 = p163 + tc;
                end
                55: begin
                        tc = f54;
                        p155 = p155 - tc;
                        p158 = p158 + tc;
                        p167 = p167 + tc;
                end
                56: begin
                        tc = f55;
                        p155 = p155 - tc;
                        p167 = p167 + tc;
                end
                57: begin
                        tc = f56;
                        p168 = p168 - tc;
                        p166 = p166 + tc;
                end
                58: begin
                        tc = f57;
                        p162 = p162 - tc;
                        p156 = p156 + tc;
                end
                59: begin
                        tc = f58;
                        p169 = p169 - tc;
                        p168 = p168 + tc;
                end
                60: begin
                        tc = f59;
                        p167 = p167 - tc;
                        p155 = p155 + tc*2;
                end
                61: begin
                        tc = f60;
                        p157 = p157 - tc;
                        p164 = p164 - tc;
                        p165 = p165 + tc;
                        p169 = p169 + tc;
                end
                62: begin
                        tc = f61;
                        p157 = p157 - tc;
                        p169 = p169 + tc;
                end
                63: begin
                        tc = f62;
                        p8 = p8 - tc;
                        p155 = p155 + tc;
                        p170 = p170 + tc;
                end
                64: begin
                        tc = f63;
                        p170 = p170 - tc;
                        p8 = p8 + tc;
                end
                65: begin
                        tc = f64;
                        p172 = p172 - tc;
                        p171 = p171 + tc;
                end
                66: begin
                        tc = f65;
                        p173 = p173 - tc;
                        p172 = p172 + tc;
                end
                67: begin
                        tc = f66;
                        p9 = p9 - tc;
                        p156 = p156 + tc;
                        p174 = p174 + tc;
                end
                68: begin
                        tc = f67;
                        p174 = p174 - tc;
                        p9 = p9 + tc;
                end
                69: begin
                        tc = f68;
                        p176 = p176 - tc;
                        p175 = p175 + tc;
                end
                70: begin
                        tc = f69;
                        p177 = p177 - tc;
                        p176 = p176 + tc;
                end
                71: begin
                        tc = f70;
                        p171 = p171 - tc;
                        p175 = p175 - tc;
                        p2 = p2 + tc;
                end
                72: begin
                        tc = f71;
                        p157 = p157 - tc;
                        p173 = p173 + tc;
                        p177 = p177 + tc;
                end
                73: begin
                        tc = f72;
                        p158 = p158 - tc;
                        p10 = p10 + tc;
                end
                74: begin
                        tc = f73;
                        p10 = p10 - tc;
                end
                75: begin
                        tc = f74;
                        p178 = p178 - tc;
                        p159 = p159 + tc;
                end
                76: begin
                        tc = f75;
                        p3 = p3 - tc;
                        p178 = p178 + tc;
                end
                77: begin
                        tc = f76;
                        p185 = p185 - tc;
                        p181 = p181 + tc;
                end
                78: begin
                        tc = f77;
                        p179 = p179 - tc;
                end
                79: begin
                        tc = f78;
                        p183 = p183 - tc;
                        p185 = p185 + tc;
                end
                80: begin
                        tc = f79;
                        p180 = p180 - tc*2;
                        p186 = p186 + tc;
                end
                81: begin
                        tc = f80;
                        p187 = p187 - tc;
                        p184 = p184 + tc;
                end
                82: begin
                        tc = f81;
                        p180 = p180 - tc;
                        p189 = p189 - tc;
                        p188 = p188 + tc;
                end
                83: begin
                        tc = f82;
                        p190 = p190 - tc;
                        p187 = p187 + tc;
                end
                84: begin
                        tc = f83;
                        p179 = p179 - tc;
                        p182 = p182 + tc;
                        p191 = p191 + tc;
                end
                85: begin
                        tc = f84;
                        p179 = p179 - tc;
                        p191 = p191 + tc;
                end
                86: begin
                        tc = f85;
                        p192 = p192 - tc;
                        p190 = p190 + tc;
                end
                87: begin
                        tc = f86;
                        p186 = p186 - tc;
                        p180 = p180 + tc;
                end
                88: begin
                        tc = f87;
                        p193 = p193 - tc;
                        p192 = p192 + tc;
                end
                89: begin
                        tc = f88;
                        p191 = p191 - tc;
                        p179 = p179 + tc*2;
                end
                90: begin
                        tc = f89;
                        p181 = p181 - tc;
                        p188 = p188 - tc;
                        p189 = p189 + tc;
                        p193 = p193 + tc;
                end
                91: begin
                        tc = f90;
                        p181 = p181 - tc;
                        p193 = p193 + tc;
                end
                92: begin
                        tc = f91;
                        p11 = p11 - tc;
                        p179 = p179 + tc;
                        p194 = p194 + tc;
                end
                93: begin
                        tc = f92;
                        p194 = p194 - tc;
                        p11 = p11 + tc;
                end
                94: begin
                        tc = f93;
                        p196 = p196 - tc;
                        p195 = p195 + tc;
                end
                95: begin
                        tc = f94;
                        p197 = p197 - tc;
                        p196 = p196 + tc;
                end
                96: begin
                        tc = f95;
                        p12 = p12 - tc;
                        p180 = p180 + tc;
                        p198 = p198 + tc;
                end
                97: begin
                        tc = f96;
                        p198 = p198 - tc;
                        p12 = p12 + tc;
                end
                98: begin
                        tc = f97;
                        p200 = p200 - tc;
                        p199 = p199 + tc;
                end
                99: begin
                        tc = f98;
                        p201 = p201 - tc;
                        p200 = p200 + tc;
                end
                100: begin
                        tc = f99;
                        p195 = p195 - tc;
                        p199 = p199 - tc;
                        p3 = p3 + tc;
                end
                101: begin
                        tc = f100;
                        p181 = p181 - tc;
                        p197 = p197 + tc;
                        p201 = p201 + tc;
                end
                102: begin
                        tc = f101;
                        p182 = p182 - tc;
                        p13 = p13 + tc;
                end
                103: begin
                        tc = f102;
                        p13 = p13 - tc;
                end
                104: begin
                        tc = f103;
                        p202 = p202 - tc;
                        p183 = p183 + tc;
                end
                105: begin
                        tc = f104;
                        p4 = p4 - tc;
                        p202 = p202 + tc;
                end
                106: begin
                        tc = f105;
                        p204 = p204 - tc;
                        p205 = p205 + tc;
                end
                107: begin
                        tc = f106;
                        p207 = p207 - tc;
                        p206 = p206 + tc;
                end
                108: begin
                        tc = f107;
                        p10 = p10 - tc;
                        p203 = p203 + tc;
                        p208 = p208 + tc;
                end
                109: begin
                        tc = f108;
                        p208 = p208 - tc;
                        p10 = p10 + tc;
                end
                110: begin
                        tc = f109;
                        p210 = p210 - tc;
                        p209 = p209 + tc;
                end
                111: begin
                        tc = f110;
                        p211 = p211 - tc;
                        p210 = p210 + tc;
                end
                112: begin
                        tc = f111;
                        p13 = p13 - tc;
                        p204 = p204 + tc;
                        p212 = p212 + tc;
                end
                113: begin
                        tc = f112;
                        p212 = p212 - tc;
                        p13 = p13 + tc;
                end
                114: begin
                        tc = f113;
                        p214 = p214 - tc;
                        p213 = p213 + tc;
                end
                115: begin
                        tc = f114;
                        p215 = p215 - tc;
                        p214 = p214 + tc;
                end
                116: begin
                        tc = f115;
                        p209 = p209 - tc;
                        p213 = p213 - tc;
                        p4 = p4 + tc;
                end
                117: begin
                        tc = f116;
                        p206 = p206 - tc;
                        p211 = p211 + tc;
                        p215 = p215 + tc;
                end
                118: begin
                        tc = f117;
                        p205 = p205 - tc;
                        p14 = p14 + tc;
                end
                119: begin
                        tc = f118;
                        p14 = p14 - tc;
                end
                120: begin
                        tc = f119;
                        p216 = p216 - tc;
                        p207 = p207 + tc;
                end
                121: begin
                        tc = f120;
                        p5 = p5 - tc;
                        p216 = p216 + tc;
                end
                122: begin
                        tc = f121;
                        p223 = p223 - tc;
                        p219 = p219 + tc;
                end
                123: begin
                        tc = f122;
                        p217 = p217 - tc;
                end
                124: begin
                        tc = f123;
                        p221 = p221 - tc;
                        p223 = p223 + tc;
                end
                125: begin
                        tc = f124;
                        p218 = p218 - tc*2;
                        p224 = p224 + tc;
                end
                126: begin
                        tc = f125;
                        p225 = p225 - tc;
                        p222 = p222 + tc;
                end
                127: begin
                        tc = f126;
                        p218 = p218 - tc;
                        p227 = p227 - tc;
                        p226 = p226 + tc;
                end
                128: begin
                        tc = f127;
                        p228 = p228 - tc;
                        p225 = p225 + tc;
                end
                129: begin
                        tc = f128;
                        p217 = p217 - tc;
                        p220 = p220 + tc;
                        p229 = p229 + tc;
                end
                130: begin
                        tc = f129;
                        p217 = p217 - tc;
                        p229 = p229 + tc;
                end
                131: begin
                        tc = f130;
                        p230 = p230 - tc;
                        p228 = p228 + tc;
                end
                132: begin
                        tc = f131;
                        p224 = p224 - tc;
                        p218 = p218 + tc;
                end
                133: begin
                        tc = f132;
                        p231 = p231 - tc;
                        p230 = p230 + tc;
                end
                134: begin
                        tc = f133;
                        p229 = p229 - tc;
                        p217 = p217 + tc*2;
                end
                135: begin
                        tc = f134;
                        p219 = p219 - tc;
                        p226 = p226 - tc;
                        p227 = p227 + tc;
                        p231 = p231 + tc;
                end
                136: begin
                        tc = f135;
                        p219 = p219 - tc;
                        p231 = p231 + tc;
                end
                137: begin
                        tc = f136;
                        p15 = p15 - tc;
                        p217 = p217 + tc;
                        p232 = p232 + tc;
                end
                138: begin
                        tc = f137;
                        p232 = p232 - tc;
                        p15 = p15 + tc;
                end
                139: begin
                        tc = f138;
                        p234 = p234 - tc;
                        p233 = p233 + tc;
                end
                140: begin
                        tc = f139;
                        p235 = p235 - tc;
                        p234 = p234 + tc;
                end
                141: begin
                        tc = f140;
                        p16 = p16 - tc;
                        p218 = p218 + tc;
                        p236 = p236 + tc;
                end
                142: begin
                        tc = f141;
                        p236 = p236 - tc;
                        p16 = p16 + tc;
                end
                143: begin
                        tc = f142;
                        p238 = p238 - tc;
                        p237 = p237 + tc;
                end
                144: begin
                        tc = f143;
                        p239 = p239 - tc;
                        p238 = p238 + tc;
                end
                145: begin
                        tc = f144;
                        p233 = p233 - tc;
                        p237 = p237 - tc;
                        p5 = p5 + tc;
                end
                146: begin
                        tc = f145;
                        p219 = p219 - tc;
                        p235 = p235 + tc;
                        p239 = p239 + tc;
                end
                147: begin
                        tc = f146;
                        p220 = p220 - tc;
                        p17 = p17 + tc;
                end
                148: begin
                        tc = f147;
                        p17 = p17 - tc;
                end
                149: begin
                        tc = f148;
                        p240 = p240 - tc;
                        p221 = p221 + tc;
                end
                150: begin
                        tc = f149;
                        p6 = p6 - tc;
                        p240 = p240 + tc;
                end
                151: begin
                        tc = f150;
                        p242 = p242 - tc;
                        p243 = p243 + tc;
                end
                152: begin
                        tc = f151;
                        p245 = p245 - tc;
                        p244 = p244 + tc;
                end
                153: begin
                        tc = f152;
                        p14 = p14 - tc;
                        p241 = p241 + tc;
                        p246 = p246 + tc;
                end
                154: begin
                        tc = f153;
                        p246 = p246 - tc;
                        p14 = p14 + tc;
                end
                155: begin
                        tc = f154;
                        p248 = p248 - tc;
                        p247 = p247 + tc;
                end
                156: begin
                        tc = f155;
                        p249 = p249 - tc;
                        p248 = p248 + tc;
                end
                157: begin
                        tc = f156;
                        p17 = p17 - tc;
                        p242 = p242 + tc;
                        p250 = p250 + tc;
                end
                158: begin
                        tc = f157;
                        p250 = p250 - tc;
                        p17 = p17 + tc;
                end
                159: begin
                        tc = f158;
                        p252 = p252 - tc;
                        p251 = p251 + tc;
                end
                160: begin
                        tc = f159;
                        p253 = p253 - tc;
                        p252 = p252 + tc;
                end
                161: begin
                        tc = f160;
                        p247 = p247 - tc;
                        p251 = p251 - tc;
                        p6 = p6 + tc;
                end
                162: begin
                        tc = f161;
                        p244 = p244 - tc;
                        p249 = p249 + tc;
                        p253 = p253 + tc;
                end
                163: begin
                        tc = f162;
                        p243 = p243 - tc;
                        p18 = p18 + tc;
                end
                164: begin
                        tc = f163;
                        p18 = p18 - tc;
                end
                165: begin
                        tc = f164;
                        p254 = p254 - tc;
                        p245 = p245 + tc;
                end
                166: begin
                        tc = f165;
                        p7 = p7 - tc;
                        p254 = p254 + tc;
                end
                167: begin
                        tc = f166;
                        p261 = p261 - tc;
                        p257 = p257 + tc;
                end
                168: begin
                        tc = f167;
                        p255 = p255 - tc;
                end
                169: begin
                        tc = f168;
                        p259 = p259 - tc;
                        p261 = p261 + tc;
                end
                170: begin
                        tc = f169;
                        p256 = p256 - tc*2;
                        p262 = p262 + tc;
                end
                171: begin
                        tc = f170;
                        p263 = p263 - tc;
                        p260 = p260 + tc;
                end
                172: begin
                        tc = f171;
                        p256 = p256 - tc;
                        p265 = p265 - tc;
                        p264 = p264 + tc;
                end
                173: begin
                        tc = f172;
                        p266 = p266 - tc;
                        p263 = p263 + tc;
                end
                174: begin
                        tc = f173;
                        p255 = p255 - tc;
                        p258 = p258 + tc;
                        p267 = p267 + tc;
                end
                175: begin
                        tc = f174;
                        p255 = p255 - tc;
                        p267 = p267 + tc;
                end
                176: begin
                        tc = f175;
                        p268 = p268 - tc;
                        p266 = p266 + tc;
                end
                177: begin
                        tc = f176;
                        p262 = p262 - tc;
                        p256 = p256 + tc;
                end
                178: begin
                        tc = f177;
                        p269 = p269 - tc;
                        p268 = p268 + tc;
                end
                179: begin
                        tc = f178;
                        p267 = p267 - tc;
                        p255 = p255 + tc*2;
                end
                180: begin
                        tc = f179;
                        p257 = p257 - tc;
                        p264 = p264 - tc;
                        p265 = p265 + tc;
                        p269 = p269 + tc;
                end
                181: begin
                        tc = f180;
                        p257 = p257 - tc;
                        p269 = p269 + tc;
                end
                182: begin
                        tc = f181;
                        p25 = p25 - tc;
                        p255 = p255 + tc;
                        p270 = p270 + tc;
                end
                183: begin
                        tc = f182;
                        p270 = p270 - tc;
                        p25 = p25 + tc;
                end
                184: begin
                        tc = f183;
                        p272 = p272 - tc;
                        p271 = p271 + tc;
                end
                185: begin
                        tc = f184;
                        p273 = p273 - tc;
                        p272 = p272 + tc;
                end
                186: begin
                        tc = f185;
                        p26 = p26 - tc;
                        p256 = p256 + tc;
                        p274 = p274 + tc;
                end
                187: begin
                        tc = f186;
                        p274 = p274 - tc;
                        p26 = p26 + tc;
                end
                188: begin
                        tc = f187;
                        p276 = p276 - tc;
                        p275 = p275 + tc;
                end
                189: begin
                        tc = f188;
                        p277 = p277 - tc;
                        p276 = p276 + tc;
                end
                190: begin
                        tc = f189;
                        p271 = p271 - tc;
                        p275 = p275 - tc;
                        p19 = p19 + tc;
                end
                191: begin
                        tc = f190;
                        p257 = p257 - tc;
                        p273 = p273 + tc;
                        p277 = p277 + tc;
                end
                192: begin
                        tc = f191;
                        p258 = p258 - tc;
                        p27 = p27 + tc;
                end
                193: begin
                        tc = f192;
                        p27 = p27 - tc;
                end
                194: begin
                        tc = f193;
                        p278 = p278 - tc;
                        p259 = p259 + tc;
                end
                195: begin
                        tc = f194;
                        p20 = p20 - tc;
                        p278 = p278 + tc;
                end
                196: begin
                        tc = f195;
                        p285 = p285 - tc;
                        p281 = p281 + tc;
                end
                197: begin
                        tc = f196;
                        p279 = p279 - tc;
                end
                198: begin
                        tc = f197;
                        p283 = p283 - tc;
                        p285 = p285 + tc;
                end
                199: begin
                        tc = f198;
                        p280 = p280 - tc*2;
                        p286 = p286 + tc;
                end
                200: begin
                        tc = f199;
                        p287 = p287 - tc;
                        p284 = p284 + tc;
                end
                201: begin
                        tc = f200;
                        p280 = p280 - tc;
                        p289 = p289 - tc;
                        p288 = p288 + tc;
                end
                202: begin
                        tc = f201;
                        p290 = p290 - tc;
                        p287 = p287 + tc;
                end
                203: begin
                        tc = f202;
                        p279 = p279 - tc;
                        p282 = p282 + tc;
                        p291 = p291 + tc;
                end
                204: begin
                        tc = f203;
                        p279 = p279 - tc;
                        p291 = p291 + tc;
                end
                205: begin
                        tc = f204;
                        p292 = p292 - tc;
                        p290 = p290 + tc;
                end
                206: begin
                        tc = f205;
                        p286 = p286 - tc;
                        p280 = p280 + tc;
                end
                207: begin
                        tc = f206;
                        p293 = p293 - tc;
                        p292 = p292 + tc;
                end
                208: begin
                        tc = f207;
                        p291 = p291 - tc;
                        p279 = p279 + tc*2;
                end
                209: begin
                        tc = f208;
                        p281 = p281 - tc;
                        p288 = p288 - tc;
                        p289 = p289 + tc;
                        p293 = p293 + tc;
                end
                210: begin
                        tc = f209;
                        p281 = p281 - tc;
                        p293 = p293 + tc;
                end
                211: begin
                        tc = f210;
                        p28 = p28 - tc;
                        p279 = p279 + tc;
                        p294 = p294 + tc;
                end
                212: begin
                        tc = f211;
                        p294 = p294 - tc;
                        p28 = p28 + tc;
                end
                213: begin
                        tc = f212;
                        p296 = p296 - tc;
                        p295 = p295 + tc;
                end
                214: begin
                        tc = f213;
                        p297 = p297 - tc;
                        p296 = p296 + tc;
                end
                215: begin
                        tc = f214;
                        p29 = p29 - tc;
                        p280 = p280 + tc;
                        p298 = p298 + tc;
                end
                216: begin
                        tc = f215;
                        p298 = p298 - tc;
                        p29 = p29 + tc;
                end
                217: begin
                        tc = f216;
                        p300 = p300 - tc;
                        p299 = p299 + tc;
                end
                218: begin
                        tc = f217;
                        p301 = p301 - tc;
                        p300 = p300 + tc;
                end
                219: begin
                        tc = f218;
                        p295 = p295 - tc;
                        p299 = p299 - tc;
                        p20 = p20 + tc;
                end
                220: begin
                        tc = f219;
                        p281 = p281 - tc;
                        p297 = p297 + tc;
                        p301 = p301 + tc;
                end
                221: begin
                        tc = f220;
                        p282 = p282 - tc;
                        p30 = p30 + tc;
                end
                222: begin
                        tc = f221;
                        p30 = p30 - tc;
                end
                223: begin
                        tc = f222;
                        p302 = p302 - tc;
                        p283 = p283 + tc;
                end
                224: begin
                        tc = f223;
                        p21 = p21 - tc;
                        p302 = p302 + tc;
                end
                225: begin
                        tc = f224;
                        p304 = p304 - tc;
                        p305 = p305 + tc;
                end
                226: begin
                        tc = f225;
                        p307 = p307 - tc;
                        p306 = p306 + tc;
                end
                227: begin
                        tc = f226;
                        p27 = p27 - tc;
                        p303 = p303 + tc;
                        p308 = p308 + tc;
                end
                228: begin
                        tc = f227;
                        p308 = p308 - tc;
                        p27 = p27 + tc;
                end
                229: begin
                        tc = f228;
                        p310 = p310 - tc;
                        p309 = p309 + tc;
                end
                230: begin
                        tc = f229;
                        p311 = p311 - tc;
                        p310 = p310 + tc;
                end
                231: begin
                        tc = f230;
                        p30 = p30 - tc;
                        p304 = p304 + tc;
                        p312 = p312 + tc;
                end
                232: begin
                        tc = f231;
                        p312 = p312 - tc;
                        p30 = p30 + tc;
                end
                233: begin
                        tc = f232;
                        p314 = p314 - tc;
                        p313 = p313 + tc;
                end
                234: begin
                        tc = f233;
                        p315 = p315 - tc;
                        p314 = p314 + tc;
                end
                235: begin
                        tc = f234;
                        p309 = p309 - tc;
                        p313 = p313 - tc;
                        p21 = p21 + tc;
                end
                236: begin
                        tc = f235;
                        p306 = p306 - tc;
                        p311 = p311 + tc;
                        p315 = p315 + tc;
                end
                237: begin
                        tc = f236;
                        p305 = p305 - tc;
                        p31 = p31 + tc;
                end
                238: begin
                        tc = f237;
                        p31 = p31 - tc;
                end
                239: begin
                        tc = f238;
                        p316 = p316 - tc;
                        p307 = p307 + tc;
                end
                240: begin
                        tc = f239;
                        p22 = p22 - tc;
                        p316 = p316 + tc;
                end
                241: begin
                        tc = f240;
                        p323 = p323 - tc;
                        p319 = p319 + tc;
                end
                242: begin
                        tc = f241;
                        p317 = p317 - tc;
                end
                243: begin
                        tc = f242;
                        p321 = p321 - tc;
                        p323 = p323 + tc;
                end
                244: begin
                        tc = f243;
                        p318 = p318 - tc*2;
                        p324 = p324 + tc;
                end
                245: begin
                        tc = f244;
                        p325 = p325 - tc;
                        p322 = p322 + tc;
                end
                246: begin
                        tc = f245;
                        p318 = p318 - tc;
                        p327 = p327 - tc;
                        p326 = p326 + tc;
                end
                247: begin
                        tc = f246;
                        p328 = p328 - tc;
                        p325 = p325 + tc;
                end
                248: begin
                        tc = f247;
                        p317 = p317 - tc;
                        p320 = p320 + tc;
                        p329 = p329 + tc;
                end
                249: begin
                        tc = f248;
                        p317 = p317 - tc;
                        p329 = p329 + tc;
                end
                250: begin
                        tc = f249;
                        p330 = p330 - tc;
                        p328 = p328 + tc;
                end
                251: begin
                        tc = f250;
                        p324 = p324 - tc;
                        p318 = p318 + tc;
                end
                252: begin
                        tc = f251;
                        p331 = p331 - tc;
                        p330 = p330 + tc;
                end
                253: begin
                        tc = f252;
                        p329 = p329 - tc;
                        p317 = p317 + tc*2;
                end
                254: begin
                        tc = f253;
                        p319 = p319 - tc;
                        p326 = p326 - tc;
                        p327 = p327 + tc;
                        p331 = p331 + tc;
                end
                255: begin
                        tc = f254;
                        p319 = p319 - tc;
                        p331 = p331 + tc;
                end
                256: begin
                        tc = f255;
                        p32 = p32 - tc;
                        p317 = p317 + tc;
                        p332 = p332 + tc;
                end
                257: begin
                        tc = f256;
                        p332 = p332 - tc;
                        p32 = p32 + tc;
                end
                258: begin
                        tc = f257;
                        p334 = p334 - tc;
                        p333 = p333 + tc;
                end
                259: begin
                        tc = f258;
                        p335 = p335 - tc;
                        p334 = p334 + tc;
                end
                260: begin
                        tc = f259;
                        p33 = p33 - tc;
                        p318 = p318 + tc;
                        p336 = p336 + tc;
                end
                261: begin
                        tc = f260;
                        p336 = p336 - tc;
                        p33 = p33 + tc;
                end
                262: begin
                        tc = f261;
                        p338 = p338 - tc;
                        p337 = p337 + tc;
                end
                263: begin
                        tc = f262;
                        p339 = p339 - tc;
                        p338 = p338 + tc;
                end
                264: begin
                        tc = f263;
                        p333 = p333 - tc;
                        p337 = p337 - tc;
                        p22 = p22 + tc;
                end
                265: begin
                        tc = f264;
                        p319 = p319 - tc;
                        p335 = p335 + tc;
                        p339 = p339 + tc;
                end
                266: begin
                        tc = f265;
                        p320 = p320 - tc;
                        p34 = p34 + tc;
                end
                267: begin
                        tc = f266;
                        p34 = p34 - tc;
                end
                268: begin
                        tc = f267;
                        p340 = p340 - tc;
                        p321 = p321 + tc;
                end
                269: begin
                        tc = f268;
                        p23 = p23 - tc;
                        p340 = p340 + tc;
                end
                270: begin
                        tc = f269;
                        p342 = p342 - tc;
                        p343 = p343 + tc;
                end
                271: begin
                        tc = f270;
                        p345 = p345 - tc;
                        p344 = p344 + tc;
                end
                272: begin
                        tc = f271;
                        p31 = p31 - tc;
                        p341 = p341 + tc;
                        p346 = p346 + tc;
                end
                273: begin
                        tc = f272;
                        p346 = p346 - tc;
                        p31 = p31 + tc;
                end
                274: begin
                        tc = f273;
                        p348 = p348 - tc;
                        p347 = p347 + tc;
                end
                275: begin
                        tc = f274;
                        p349 = p349 - tc;
                        p348 = p348 + tc;
                end
                276: begin
                        tc = f275;
                        p34 = p34 - tc;
                        p342 = p342 + tc;
                        p350 = p350 + tc;
                end
                277: begin
                        tc = f276;
                        p350 = p350 - tc;
                        p34 = p34 + tc;
                end
                278: begin
                        tc = f277;
                        p352 = p352 - tc;
                        p351 = p351 + tc;
                end
                279: begin
                        tc = f278;
                        p353 = p353 - tc;
                        p352 = p352 + tc;
                end
                280: begin
                        tc = f279;
                        p347 = p347 - tc;
                        p351 = p351 - tc;
                        p23 = p23 + tc;
                end
                281: begin
                        tc = f280;
                        p344 = p344 - tc;
                        p349 = p349 + tc;
                        p353 = p353 + tc;
                end
                282: begin
                        tc = f281;
                        p343 = p343 - tc;
                        p35 = p35 + tc;
                end
                283: begin
                        tc = f282;
                        p35 = p35 - tc;
                end
                284: begin
                        tc = f283;
                        p354 = p354 - tc;
                        p345 = p345 + tc;
                end
                285: begin
                        tc = f284;
                        p24 = p24 - tc;
                        p354 = p354 + tc;
                end
                286: begin
                        tc = f285;
                        p361 = p361 - tc;
                        p357 = p357 + tc;
                end
                287: begin
                        tc = f286;
                        p355 = p355 - tc;
                end
                288: begin
                        tc = f287;
                        p359 = p359 - tc;
                        p361 = p361 + tc;
                end
                289: begin
                        tc = f288;
                        p356 = p356 - tc*2;
                        p362 = p362 + tc;
                end
                290: begin
                        tc = f289;
                        p363 = p363 - tc;
                        p360 = p360 + tc;
                end
                291: begin
                        tc = f290;
                        p356 = p356 - tc;
                        p365 = p365 - tc;
                        p364 = p364 + tc;
                end
                292: begin
                        tc = f291;
                        p366 = p366 - tc;
                        p363 = p363 + tc;
                end
                293: begin
                        tc = f292;
                        p355 = p355 - tc;
                        p358 = p358 + tc;
                        p367 = p367 + tc;
                end
                294: begin
                        tc = f293;
                        p355 = p355 - tc;
                        p367 = p367 + tc;
                end
                295: begin
                        tc = f294;
                        p368 = p368 - tc;
                        p366 = p366 + tc;
                end
                296: begin
                        tc = f295;
                        p362 = p362 - tc;
                        p356 = p356 + tc;
                end
                297: begin
                        tc = f296;
                        p369 = p369 - tc;
                        p368 = p368 + tc;
                end
                298: begin
                        tc = f297;
                        p367 = p367 - tc;
                        p355 = p355 + tc*2;
                end
                299: begin
                        tc = f298;
                        p357 = p357 - tc;
                        p364 = p364 - tc;
                        p365 = p365 + tc;
                        p369 = p369 + tc;
                end
                300: begin
                        tc = f299;
                        p357 = p357 - tc;
                        p369 = p369 + tc;
                end
                301: begin
                        tc = f300;
                        p42 = p42 - tc;
                        p355 = p355 + tc;
                        p370 = p370 + tc;
                end
                302: begin
                        tc = f301;
                        p370 = p370 - tc;
                        p42 = p42 + tc;
                end
                303: begin
                        tc = f302;
                        p372 = p372 - tc;
                        p371 = p371 + tc;
                end
                304: begin
                        tc = f303;
                        p373 = p373 - tc;
                        p372 = p372 + tc;
                end
                305: begin
                        tc = f304;
                        p43 = p43 - tc;
                        p356 = p356 + tc;
                        p374 = p374 + tc;
                end
                306: begin
                        tc = f305;
                        p374 = p374 - tc;
                        p43 = p43 + tc;
                end
                307: begin
                        tc = f306;
                        p376 = p376 - tc;
                        p375 = p375 + tc;
                end
                308: begin
                        tc = f307;
                        p377 = p377 - tc;
                        p376 = p376 + tc;
                end
                309: begin
                        tc = f308;
                        p371 = p371 - tc;
                        p375 = p375 - tc;
                        p36 = p36 + tc;
                end
                310: begin
                        tc = f309;
                        p357 = p357 - tc;
                        p373 = p373 + tc;
                        p377 = p377 + tc;
                end
                311: begin
                        tc = f310;
                        p358 = p358 - tc;
                        p44 = p44 + tc;
                end
                312: begin
                        tc = f311;
                        p44 = p44 - tc;
                end
                313: begin
                        tc = f312;
                        p378 = p378 - tc;
                        p359 = p359 + tc;
                end
                314: begin
                        tc = f313;
                        p37 = p37 - tc;
                        p378 = p378 + tc;
                end
                315: begin
                        tc = f314;
                        p385 = p385 - tc;
                        p381 = p381 + tc;
                end
                316: begin
                        tc = f315;
                        p379 = p379 - tc;
                end
                317: begin
                        tc = f316;
                        p383 = p383 - tc;
                        p385 = p385 + tc;
                end
                318: begin
                        tc = f317;
                        p380 = p380 - tc*2;
                        p386 = p386 + tc;
                end
                319: begin
                        tc = f318;
                        p387 = p387 - tc;
                        p384 = p384 + tc;
                end
                320: begin
                        tc = f319;
                        p380 = p380 - tc;
                        p389 = p389 - tc;
                        p388 = p388 + tc;
                end
                321: begin
                        tc = f320;
                        p390 = p390 - tc;
                        p387 = p387 + tc;
                end
                322: begin
                        tc = f321;
                        p379 = p379 - tc;
                        p382 = p382 + tc;
                        p391 = p391 + tc;
                end
                323: begin
                        tc = f322;
                        p379 = p379 - tc;
                        p391 = p391 + tc;
                end
                324: begin
                        tc = f323;
                        p392 = p392 - tc;
                        p390 = p390 + tc;
                end
                325: begin
                        tc = f324;
                        p386 = p386 - tc;
                        p380 = p380 + tc;
                end
                326: begin
                        tc = f325;
                        p393 = p393 - tc;
                        p392 = p392 + tc;
                end
                327: begin
                        tc = f326;
                        p391 = p391 - tc;
                        p379 = p379 + tc*2;
                end
                328: begin
                        tc = f327;
                        p381 = p381 - tc;
                        p388 = p388 - tc;
                        p389 = p389 + tc;
                        p393 = p393 + tc;
                end
                329: begin
                        tc = f328;
                        p381 = p381 - tc;
                        p393 = p393 + tc;
                end
                330: begin
                        tc = f329;
                        p45 = p45 - tc;
                        p379 = p379 + tc;
                        p394 = p394 + tc;
                end
                331: begin
                        tc = f330;
                        p394 = p394 - tc;
                        p45 = p45 + tc;
                end
                332: begin
                        tc = f331;
                        p396 = p396 - tc;
                        p395 = p395 + tc;
                end
                333: begin
                        tc = f332;
                        p397 = p397 - tc;
                        p396 = p396 + tc;
                end
                334: begin
                        tc = f333;
                        p46 = p46 - tc;
                        p380 = p380 + tc;
                        p398 = p398 + tc;
                end
                335: begin
                        tc = f334;
                        p398 = p398 - tc;
                        p46 = p46 + tc;
                end
                336: begin
                        tc = f335;
                        p400 = p400 - tc;
                        p399 = p399 + tc;
                end
                337: begin
                        tc = f336;
                        p401 = p401 - tc;
                        p400 = p400 + tc;
                end
                338: begin
                        tc = f337;
                        p395 = p395 - tc;
                        p399 = p399 - tc;
                        p37 = p37 + tc;
                end
                339: begin
                        tc = f338;
                        p381 = p381 - tc;
                        p397 = p397 + tc;
                        p401 = p401 + tc;
                end
                340: begin
                        tc = f339;
                        p382 = p382 - tc;
                        p47 = p47 + tc;
                end
                341: begin
                        tc = f340;
                        p47 = p47 - tc;
                end
                342: begin
                        tc = f341;
                        p402 = p402 - tc;
                        p383 = p383 + tc;
                end
                343: begin
                        tc = f342;
                        p38 = p38 - tc;
                        p402 = p402 + tc;
                end
                344: begin
                        tc = f343;
                        p404 = p404 - tc;
                        p405 = p405 + tc;
                end
                345: begin
                        tc = f344;
                        p407 = p407 - tc;
                        p406 = p406 + tc;
                end
                346: begin
                        tc = f345;
                        p44 = p44 - tc;
                        p403 = p403 + tc;
                        p408 = p408 + tc;
                end
                347: begin
                        tc = f346;
                        p408 = p408 - tc;
                        p44 = p44 + tc;
                end
                348: begin
                        tc = f347;
                        p410 = p410 - tc;
                        p409 = p409 + tc;
                end
                349: begin
                        tc = f348;
                        p411 = p411 - tc;
                        p410 = p410 + tc;
                end
                350: begin
                        tc = f349;
                        p47 = p47 - tc;
                        p404 = p404 + tc;
                        p412 = p412 + tc;
                end
                351: begin
                        tc = f350;
                        p412 = p412 - tc;
                        p47 = p47 + tc;
                end
                352: begin
                        tc = f351;
                        p414 = p414 - tc;
                        p413 = p413 + tc;
                end
                353: begin
                        tc = f352;
                        p415 = p415 - tc;
                        p414 = p414 + tc;
                end
                354: begin
                        tc = f353;
                        p409 = p409 - tc;
                        p413 = p413 - tc;
                        p38 = p38 + tc;
                end
                355: begin
                        tc = f354;
                        p406 = p406 - tc;
                        p411 = p411 + tc;
                        p415 = p415 + tc;
                end
                356: begin
                        tc = f355;
                        p405 = p405 - tc;
                        p48 = p48 + tc;
                end
                357: begin
                        tc = f356;
                        p48 = p48 - tc;
                end
                358: begin
                        tc = f357;
                        p416 = p416 - tc;
                        p407 = p407 + tc;
                end
                359: begin
                        tc = f358;
                        p39 = p39 - tc;
                        p416 = p416 + tc;
                end
                360: begin
                        tc = f359;
                        p423 = p423 - tc;
                        p419 = p419 + tc;
                end
                361: begin
                        tc = f360;
                        p417 = p417 - tc;
                end
                362: begin
                        tc = f361;
                        p421 = p421 - tc;
                        p423 = p423 + tc;
                end
                363: begin
                        tc = f362;
                        p418 = p418 - tc*2;
                        p424 = p424 + tc;
                end
                364: begin
                        tc = f363;
                        p425 = p425 - tc;
                        p422 = p422 + tc;
                end
                365: begin
                        tc = f364;
                        p418 = p418 - tc;
                        p427 = p427 - tc;
                        p426 = p426 + tc;
                end
                366: begin
                        tc = f365;
                        p428 = p428 - tc;
                        p425 = p425 + tc;
                end
                367: begin
                        tc = f366;
                        p417 = p417 - tc;
                        p420 = p420 + tc;
                        p429 = p429 + tc;
                end
                368: begin
                        tc = f367;
                        p417 = p417 - tc;
                        p429 = p429 + tc;
                end
                369: begin
                        tc = f368;
                        p430 = p430 - tc;
                        p428 = p428 + tc;
                end
                370: begin
                        tc = f369;
                        p424 = p424 - tc;
                        p418 = p418 + tc;
                end
                371: begin
                        tc = f370;
                        p431 = p431 - tc;
                        p430 = p430 + tc;
                end
                372: begin
                        tc = f371;
                        p429 = p429 - tc;
                        p417 = p417 + tc*2;
                end
                373: begin
                        tc = f372;
                        p419 = p419 - tc;
                        p426 = p426 - tc;
                        p427 = p427 + tc;
                        p431 = p431 + tc;
                end
                374: begin
                        tc = f373;
                        p419 = p419 - tc;
                        p431 = p431 + tc;
                end
                375: begin
                        tc = f374;
                        p49 = p49 - tc;
                        p417 = p417 + tc;
                        p432 = p432 + tc;
                end
                376: begin
                        tc = f375;
                        p432 = p432 - tc;
                        p49 = p49 + tc;
                end
                377: begin
                        tc = f376;
                        p434 = p434 - tc;
                        p433 = p433 + tc;
                end
                378: begin
                        tc = f377;
                        p435 = p435 - tc;
                        p434 = p434 + tc;
                end
                379: begin
                        tc = f378;
                        p50 = p50 - tc;
                        p418 = p418 + tc;
                        p436 = p436 + tc;
                end
                380: begin
                        tc = f379;
                        p436 = p436 - tc;
                        p50 = p50 + tc;
                end
                381: begin
                        tc = f380;
                        p438 = p438 - tc;
                        p437 = p437 + tc;
                end
                382: begin
                        tc = f381;
                        p439 = p439 - tc;
                        p438 = p438 + tc;
                end
                383: begin
                        tc = f382;
                        p433 = p433 - tc;
                        p437 = p437 - tc;
                        p39 = p39 + tc;
                end
                384: begin
                        tc = f383;
                        p419 = p419 - tc;
                        p435 = p435 + tc;
                        p439 = p439 + tc;
                end
                385: begin
                        tc = f384;
                        p420 = p420 - tc;
                        p51 = p51 + tc;
                end
                386: begin
                        tc = f385;
                        p51 = p51 - tc;
                end
                387: begin
                        tc = f386;
                        p440 = p440 - tc;
                        p421 = p421 + tc;
                end
                388: begin
                        tc = f387;
                        p40 = p40 - tc;
                        p440 = p440 + tc;
                end
                389: begin
                        tc = f388;
                        p442 = p442 - tc;
                        p443 = p443 + tc;
                end
                390: begin
                        tc = f389;
                        p445 = p445 - tc;
                        p444 = p444 + tc;
                end
                391: begin
                        tc = f390;
                        p48 = p48 - tc;
                        p441 = p441 + tc;
                        p446 = p446 + tc;
                end
                392: begin
                        tc = f391;
                        p446 = p446 - tc;
                        p48 = p48 + tc;
                end
                393: begin
                        tc = f392;
                        p448 = p448 - tc;
                        p447 = p447 + tc;
                end
                394: begin
                        tc = f393;
                        p449 = p449 - tc;
                        p448 = p448 + tc;
                end
                395: begin
                        tc = f394;
                        p51 = p51 - tc;
                        p442 = p442 + tc;
                        p450 = p450 + tc;
                end
                396: begin
                        tc = f395;
                        p450 = p450 - tc;
                        p51 = p51 + tc;
                end
                397: begin
                        tc = f396;
                        p452 = p452 - tc;
                        p451 = p451 + tc;
                end
                398: begin
                        tc = f397;
                        p453 = p453 - tc;
                        p452 = p452 + tc;
                end
                399: begin
                        tc = f398;
                        p447 = p447 - tc;
                        p451 = p451 - tc;
                        p40 = p40 + tc;
                end
                400: begin
                        tc = f399;
                        p444 = p444 - tc;
                        p449 = p449 + tc;
                        p453 = p453 + tc;
                end
                401: begin
                        tc = f400;
                        p443 = p443 - tc;
                        p52 = p52 + tc;
                end
                402: begin
                        tc = f401;
                        p52 = p52 - tc;
                end
                403: begin
                        tc = f402;
                        p454 = p454 - tc;
                        p445 = p445 + tc;
                end
                404: begin
                        tc = f403;
                        p41 = p41 - tc;
                        p454 = p454 + tc;
                end
                405: begin
                        tc = f404;
                        p461 = p461 - tc;
                        p457 = p457 + tc;
                end
                406: begin
                        tc = f405;
                        p455 = p455 - tc;
                end
                407: begin
                        tc = f406;
                        p459 = p459 - tc;
                        p461 = p461 + tc;
                end
                408: begin
                        tc = f407;
                        p456 = p456 - tc*2;
                        p462 = p462 + tc;
                end
                409: begin
                        tc = f408;
                        p463 = p463 - tc;
                        p460 = p460 + tc;
                end
                410: begin
                        tc = f409;
                        p456 = p456 - tc;
                        p465 = p465 - tc;
                        p464 = p464 + tc;
                end
                411: begin
                        tc = f410;
                        p466 = p466 - tc;
                        p463 = p463 + tc;
                end
                412: begin
                        tc = f411;
                        p455 = p455 - tc;
                        p458 = p458 + tc;
                        p467 = p467 + tc;
                end
                413: begin
                        tc = f412;
                        p455 = p455 - tc;
                        p467 = p467 + tc;
                end
                414: begin
                        tc = f413;
                        p468 = p468 - tc;
                        p466 = p466 + tc;
                end
                415: begin
                        tc = f414;
                        p462 = p462 - tc;
                        p456 = p456 + tc;
                end
                416: begin
                        tc = f415;
                        p469 = p469 - tc;
                        p468 = p468 + tc;
                end
                417: begin
                        tc = f416;
                        p467 = p467 - tc;
                        p455 = p455 + tc*2;
                end
                418: begin
                        tc = f417;
                        p457 = p457 - tc;
                        p464 = p464 - tc;
                        p465 = p465 + tc;
                        p469 = p469 + tc;
                end
                419: begin
                        tc = f418;
                        p457 = p457 - tc;
                        p469 = p469 + tc;
                end
                420: begin
                        tc = f419;
                        p59 = p59 - tc;
                        p455 = p455 + tc;
                        p470 = p470 + tc;
                end
                421: begin
                        tc = f420;
                        p470 = p470 - tc;
                        p59 = p59 + tc;
                end
                422: begin
                        tc = f421;
                        p472 = p472 - tc;
                        p471 = p471 + tc;
                end
                423: begin
                        tc = f422;
                        p473 = p473 - tc;
                        p472 = p472 + tc;
                end
                424: begin
                        tc = f423;
                        p60 = p60 - tc;
                        p456 = p456 + tc;
                        p474 = p474 + tc;
                end
                425: begin
                        tc = f424;
                        p474 = p474 - tc;
                        p60 = p60 + tc;
                end
                426: begin
                        tc = f425;
                        p476 = p476 - tc;
                        p475 = p475 + tc;
                end
                427: begin
                        tc = f426;
                        p477 = p477 - tc;
                        p476 = p476 + tc;
                end
                428: begin
                        tc = f427;
                        p471 = p471 - tc;
                        p475 = p475 - tc;
                        p53 = p53 + tc;
                end
                429: begin
                        tc = f428;
                        p457 = p457 - tc;
                        p473 = p473 + tc;
                        p477 = p477 + tc;
                end
                430: begin
                        tc = f429;
                        p458 = p458 - tc;
                        p61 = p61 + tc;
                end
                431: begin
                        tc = f430;
                        p61 = p61 - tc;
                end
                432: begin
                        tc = f431;
                        p478 = p478 - tc;
                        p459 = p459 + tc;
                end
                433: begin
                        tc = f432;
                        p54 = p54 - tc;
                        p478 = p478 + tc;
                end
                434: begin
                        tc = f433;
                        p485 = p485 - tc;
                        p481 = p481 + tc;
                end
                435: begin
                        tc = f434;
                        p479 = p479 - tc;
                end
                436: begin
                        tc = f435;
                        p483 = p483 - tc;
                        p485 = p485 + tc;
                end
                437: begin
                        tc = f436;
                        p480 = p480 - tc*2;
                        p486 = p486 + tc;
                end
                438: begin
                        tc = f437;
                        p487 = p487 - tc;
                        p484 = p484 + tc;
                end
                439: begin
                        tc = f438;
                        p480 = p480 - tc;
                        p489 = p489 - tc;
                        p488 = p488 + tc;
                end
                440: begin
                        tc = f439;
                        p490 = p490 - tc;
                        p487 = p487 + tc;
                end
                441: begin
                        tc = f440;
                        p479 = p479 - tc;
                        p482 = p482 + tc;
                        p491 = p491 + tc;
                end
                442: begin
                        tc = f441;
                        p479 = p479 - tc;
                        p491 = p491 + tc;
                end
                443: begin
                        tc = f442;
                        p492 = p492 - tc;
                        p490 = p490 + tc;
                end
                444: begin
                        tc = f443;
                        p486 = p486 - tc;
                        p480 = p480 + tc;
                end
                445: begin
                        tc = f444;
                        p493 = p493 - tc;
                        p492 = p492 + tc;
                end
                446: begin
                        tc = f445;
                        p491 = p491 - tc;
                        p479 = p479 + tc*2;
                end
                447: begin
                        tc = f446;
                        p481 = p481 - tc;
                        p488 = p488 - tc;
                        p489 = p489 + tc;
                        p493 = p493 + tc;
                end
                448: begin
                        tc = f447;
                        p481 = p481 - tc;
                        p493 = p493 + tc;
                end
                449: begin
                        tc = f448;
                        p62 = p62 - tc;
                        p479 = p479 + tc;
                        p494 = p494 + tc;
                end
                450: begin
                        tc = f449;
                        p494 = p494 - tc;
                        p62 = p62 + tc;
                end
                451: begin
                        tc = f450;
                        p496 = p496 - tc;
                        p495 = p495 + tc;
                end
                452: begin
                        tc = f451;
                        p497 = p497 - tc;
                        p496 = p496 + tc;
                end
                453: begin
                        tc = f452;
                        p63 = p63 - tc;
                        p480 = p480 + tc;
                        p498 = p498 + tc;
                end
                454: begin
                        tc = f453;
                        p498 = p498 - tc;
                        p63 = p63 + tc;
                end
                455: begin
                        tc = f454;
                        p500 = p500 - tc;
                        p499 = p499 + tc;
                end
                456: begin
                        tc = f455;
                        p501 = p501 - tc;
                        p500 = p500 + tc;
                end
                457: begin
                        tc = f456;
                        p495 = p495 - tc;
                        p499 = p499 - tc;
                        p54 = p54 + tc;
                end
                458: begin
                        tc = f457;
                        p481 = p481 - tc;
                        p497 = p497 + tc;
                        p501 = p501 + tc;
                end
                459: begin
                        tc = f458;
                        p482 = p482 - tc;
                        p64 = p64 + tc;
                end
                460: begin
                        tc = f459;
                        p64 = p64 - tc;
                end
                461: begin
                        tc = f460;
                        p502 = p502 - tc;
                        p483 = p483 + tc;
                end
                462: begin
                        tc = f461;
                        p55 = p55 - tc;
                        p502 = p502 + tc;
                end
                463: begin
                        tc = f462;
                        p504 = p504 - tc;
                        p505 = p505 + tc;
                end
                464: begin
                        tc = f463;
                        p507 = p507 - tc;
                        p506 = p506 + tc;
                end
                465: begin
                        tc = f464;
                        p61 = p61 - tc;
                        p503 = p503 + tc;
                        p508 = p508 + tc;
                end
                466: begin
                        tc = f465;
                        p508 = p508 - tc;
                        p61 = p61 + tc;
                end
                467: begin
                        tc = f466;
                        p510 = p510 - tc;
                        p509 = p509 + tc;
                end
                468: begin
                        tc = f467;
                        p511 = p511 - tc;
                        p510 = p510 + tc;
                end
                469: begin
                        tc = f468;
                        p64 = p64 - tc;
                        p504 = p504 + tc;
                        p512 = p512 + tc;
                end
                470: begin
                        tc = f469;
                        p512 = p512 - tc;
                        p64 = p64 + tc;
                end
                471: begin
                        tc = f470;
                        p514 = p514 - tc;
                        p513 = p513 + tc;
                end
                472: begin
                        tc = f471;
                        p515 = p515 - tc;
                        p514 = p514 + tc;
                end
                473: begin
                        tc = f472;
                        p509 = p509 - tc;
                        p513 = p513 - tc;
                        p55 = p55 + tc;
                end
                474: begin
                        tc = f473;
                        p506 = p506 - tc;
                        p511 = p511 + tc;
                        p515 = p515 + tc;
                end
                475: begin
                        tc = f474;
                        p505 = p505 - tc;
                        p65 = p65 + tc;
                end
                476: begin
                        tc = f475;
                        p65 = p65 - tc;
                end
                477: begin
                        tc = f476;
                        p516 = p516 - tc;
                        p507 = p507 + tc;
                end
                478: begin
                        tc = f477;
                        p56 = p56 - tc;
                        p516 = p516 + tc;
                end
                479: begin
                        tc = f478;
                        p523 = p523 - tc;
                        p519 = p519 + tc;
                end
                480: begin
                        tc = f479;
                        p517 = p517 - tc;
                end
                481: begin
                        tc = f480;
                        p521 = p521 - tc;
                        p523 = p523 + tc;
                end
                482: begin
                        tc = f481;
                        p518 = p518 - tc*2;
                        p524 = p524 + tc;
                end
                483: begin
                        tc = f482;
                        p525 = p525 - tc;
                        p522 = p522 + tc;
                end
                484: begin
                        tc = f483;
                        p518 = p518 - tc;
                        p527 = p527 - tc;
                        p526 = p526 + tc;
                end
                485: begin
                        tc = f484;
                        p528 = p528 - tc;
                        p525 = p525 + tc;
                end
                486: begin
                        tc = f485;
                        p517 = p517 - tc;
                        p520 = p520 + tc;
                        p529 = p529 + tc;
                end
                487: begin
                        tc = f486;
                        p517 = p517 - tc;
                        p529 = p529 + tc;
                end
                488: begin
                        tc = f487;
                        p530 = p530 - tc;
                        p528 = p528 + tc;
                end
                489: begin
                        tc = f488;
                        p524 = p524 - tc;
                        p518 = p518 + tc;
                end
                490: begin
                        tc = f489;
                        p531 = p531 - tc;
                        p530 = p530 + tc;
                end
                491: begin
                        tc = f490;
                        p529 = p529 - tc;
                        p517 = p517 + tc*2;
                end
                492: begin
                        tc = f491;
                        p519 = p519 - tc;
                        p526 = p526 - tc;
                        p527 = p527 + tc;
                        p531 = p531 + tc;
                end
                493: begin
                        tc = f492;
                        p519 = p519 - tc;
                        p531 = p531 + tc;
                end
                494: begin
                        tc = f493;
                        p66 = p66 - tc;
                        p517 = p517 + tc;
                        p532 = p532 + tc;
                end
                495: begin
                        tc = f494;
                        p532 = p532 - tc;
                        p66 = p66 + tc;
                end
                496: begin
                        tc = f495;
                        p534 = p534 - tc;
                        p533 = p533 + tc;
                end
                497: begin
                        tc = f496;
                        p535 = p535 - tc;
                        p534 = p534 + tc;
                end
                498: begin
                        tc = f497;
                        p67 = p67 - tc;
                        p518 = p518 + tc;
                        p536 = p536 + tc;
                end
                499: begin
                        tc = f498;
                        p536 = p536 - tc;
                        p67 = p67 + tc;
                end
                500: begin
                        tc = f499;
                        p538 = p538 - tc;
                        p537 = p537 + tc;
                end
                501: begin
                        tc = f500;
                        p539 = p539 - tc;
                        p538 = p538 + tc;
                end
                502: begin
                        tc = f501;
                        p533 = p533 - tc;
                        p537 = p537 - tc;
                        p56 = p56 + tc;
                end
                503: begin
                        tc = f502;
                        p519 = p519 - tc;
                        p535 = p535 + tc;
                        p539 = p539 + tc;
                end
                504: begin
                        tc = f503;
                        p520 = p520 - tc;
                        p68 = p68 + tc;
                end
                505: begin
                        tc = f504;
                        p68 = p68 - tc;
                end
                506: begin
                        tc = f505;
                        p540 = p540 - tc;
                        p521 = p521 + tc;
                end
                507: begin
                        tc = f506;
                        p57 = p57 - tc;
                        p540 = p540 + tc;
                end
                508: begin
                        tc = f507;
                        p542 = p542 - tc;
                        p543 = p543 + tc;
                end
                509: begin
                        tc = f508;
                        p545 = p545 - tc;
                        p544 = p544 + tc;
                end
                510: begin
                        tc = f509;
                        p65 = p65 - tc;
                        p541 = p541 + tc;
                        p546 = p546 + tc;
                end
                511: begin
                        tc = f510;
                        p546 = p546 - tc;
                        p65 = p65 + tc;
                end
                512: begin
                        tc = f511;
                        p548 = p548 - tc;
                        p547 = p547 + tc;
                end
                513: begin
                        tc = f512;
                        p549 = p549 - tc;
                        p548 = p548 + tc;
                end
                514: begin
                        tc = f513;
                        p68 = p68 - tc;
                        p542 = p542 + tc;
                        p550 = p550 + tc;
                end
                515: begin
                        tc = f514;
                        p550 = p550 - tc;
                        p68 = p68 + tc;
                end
                516: begin
                        tc = f515;
                        p552 = p552 - tc;
                        p551 = p551 + tc;
                end
                517: begin
                        tc = f516;
                        p553 = p553 - tc;
                        p552 = p552 + tc;
                end
                518: begin
                        tc = f517;
                        p547 = p547 - tc;
                        p551 = p551 - tc;
                        p57 = p57 + tc;
                end
                519: begin
                        tc = f518;
                        p544 = p544 - tc;
                        p549 = p549 + tc;
                        p553 = p553 + tc;
                end
                520: begin
                        tc = f519;
                        p543 = p543 - tc;
                        p69 = p69 + tc;
                end
                521: begin
                        tc = f520;
                        p69 = p69 - tc;
                end
                522: begin
                        tc = f521;
                        p554 = p554 - tc;
                        p545 = p545 + tc;
                end
                523: begin
                        tc = f522;
                        p58 = p58 - tc;
                        p554 = p554 + tc;
                end
                524: begin
                        tc = f523;
                        p561 = p561 - tc;
                        p557 = p557 + tc;
                end
                525: begin
                        tc = f524;
                        p555 = p555 - tc;
                end
                526: begin
                        tc = f525;
                        p559 = p559 - tc;
                        p561 = p561 + tc;
                end
                527: begin
                        tc = f526;
                        p556 = p556 - tc*2;
                        p562 = p562 + tc;
                end
                528: begin
                        tc = f527;
                        p563 = p563 - tc;
                        p560 = p560 + tc;
                end
                529: begin
                        tc = f528;
                        p556 = p556 - tc;
                        p565 = p565 - tc;
                        p564 = p564 + tc;
                end
                530: begin
                        tc = f529;
                        p566 = p566 - tc;
                        p563 = p563 + tc;
                end
                531: begin
                        tc = f530;
                        p555 = p555 - tc;
                        p558 = p558 + tc;
                        p567 = p567 + tc;
                end
                532: begin
                        tc = f531;
                        p555 = p555 - tc;
                        p567 = p567 + tc;
                end
                533: begin
                        tc = f532;
                        p568 = p568 - tc;
                        p566 = p566 + tc;
                end
                534: begin
                        tc = f533;
                        p562 = p562 - tc;
                        p556 = p556 + tc;
                end
                535: begin
                        tc = f534;
                        p569 = p569 - tc;
                        p568 = p568 + tc;
                end
                536: begin
                        tc = f535;
                        p567 = p567 - tc;
                        p555 = p555 + tc*2;
                end
                537: begin
                        tc = f536;
                        p557 = p557 - tc;
                        p564 = p564 - tc;
                        p565 = p565 + tc;
                        p569 = p569 + tc;
                end
                538: begin
                        tc = f537;
                        p557 = p557 - tc;
                        p569 = p569 + tc;
                end
                539: begin
                        tc = f538;
                        p76 = p76 - tc;
                        p555 = p555 + tc;
                        p570 = p570 + tc;
                end
                540: begin
                        tc = f539;
                        p570 = p570 - tc;
                        p76 = p76 + tc;
                end
                541: begin
                        tc = f540;
                        p572 = p572 - tc;
                        p571 = p571 + tc;
                end
                542: begin
                        tc = f541;
                        p573 = p573 - tc;
                        p572 = p572 + tc;
                end
                543: begin
                        tc = f542;
                        p77 = p77 - tc;
                        p556 = p556 + tc;
                        p574 = p574 + tc;
                end
                544: begin
                        tc = f543;
                        p574 = p574 - tc;
                        p77 = p77 + tc;
                end
                545: begin
                        tc = f544;
                        p576 = p576 - tc;
                        p575 = p575 + tc;
                end
                546: begin
                        tc = f545;
                        p577 = p577 - tc;
                        p576 = p576 + tc;
                end
                547: begin
                        tc = f546;
                        p571 = p571 - tc;
                        p575 = p575 - tc;
                        p70 = p70 + tc;
                end
                548: begin
                        tc = f547;
                        p557 = p557 - tc;
                        p573 = p573 + tc;
                        p577 = p577 + tc;
                end
                549: begin
                        tc = f548;
                        p558 = p558 - tc;
                        p78 = p78 + tc;
                end
                550: begin
                        tc = f549;
                        p78 = p78 - tc;
                end
                551: begin
                        tc = f550;
                        p578 = p578 - tc;
                        p559 = p559 + tc;
                end
                552: begin
                        tc = f551;
                        p71 = p71 - tc;
                        p578 = p578 + tc;
                end
                553: begin
                        tc = f552;
                        p585 = p585 - tc;
                        p581 = p581 + tc;
                end
                554: begin
                        tc = f553;
                        p579 = p579 - tc;
                end
                555: begin
                        tc = f554;
                        p583 = p583 - tc;
                        p585 = p585 + tc;
                end
                556: begin
                        tc = f555;
                        p580 = p580 - tc*2;
                        p586 = p586 + tc;
                end
                557: begin
                        tc = f556;
                        p587 = p587 - tc;
                        p584 = p584 + tc;
                end
                558: begin
                        tc = f557;
                        p580 = p580 - tc;
                        p589 = p589 - tc;
                        p588 = p588 + tc;
                end
                559: begin
                        tc = f558;
                        p590 = p590 - tc;
                        p587 = p587 + tc;
                end
                560: begin
                        tc = f559;
                        p579 = p579 - tc;
                        p582 = p582 + tc;
                        p591 = p591 + tc;
                end
                561: begin
                        tc = f560;
                        p579 = p579 - tc;
                        p591 = p591 + tc;
                end
                562: begin
                        tc = f561;
                        p592 = p592 - tc;
                        p590 = p590 + tc;
                end
                563: begin
                        tc = f562;
                        p586 = p586 - tc;
                        p580 = p580 + tc;
                end
                564: begin
                        tc = f563;
                        p593 = p593 - tc;
                        p592 = p592 + tc;
                end
                565: begin
                        tc = f564;
                        p591 = p591 - tc;
                        p579 = p579 + tc*2;
                end
                566: begin
                        tc = f565;
                        p581 = p581 - tc;
                        p588 = p588 - tc;
                        p589 = p589 + tc;
                        p593 = p593 + tc;
                end
                567: begin
                        tc = f566;
                        p581 = p581 - tc;
                        p593 = p593 + tc;
                end
                568: begin
                        tc = f567;
                        p79 = p79 - tc;
                        p579 = p579 + tc;
                        p594 = p594 + tc;
                end
                569: begin
                        tc = f568;
                        p594 = p594 - tc;
                        p79 = p79 + tc;
                end
                570: begin
                        tc = f569;
                        p596 = p596 - tc;
                        p595 = p595 + tc;
                end
                571: begin
                        tc = f570;
                        p597 = p597 - tc;
                        p596 = p596 + tc;
                end
                572: begin
                        tc = f571;
                        p80 = p80 - tc;
                        p580 = p580 + tc;
                        p598 = p598 + tc;
                end
                573: begin
                        tc = f572;
                        p598 = p598 - tc;
                        p80 = p80 + tc;
                end
                574: begin
                        tc = f573;
                        p600 = p600 - tc;
                        p599 = p599 + tc;
                end
                575: begin
                        tc = f574;
                        p601 = p601 - tc;
                        p600 = p600 + tc;
                end
                576: begin
                        tc = f575;
                        p595 = p595 - tc;
                        p599 = p599 - tc;
                        p71 = p71 + tc;
                end
                577: begin
                        tc = f576;
                        p581 = p581 - tc;
                        p597 = p597 + tc;
                        p601 = p601 + tc;
                end
                578: begin
                        tc = f577;
                        p582 = p582 - tc;
                        p81 = p81 + tc;
                end
                579: begin
                        tc = f578;
                        p81 = p81 - tc;
                end
                580: begin
                        tc = f579;
                        p602 = p602 - tc;
                        p583 = p583 + tc;
                end
                581: begin
                        tc = f580;
                        p72 = p72 - tc;
                        p602 = p602 + tc;
                end
                582: begin
                        tc = f581;
                        p604 = p604 - tc;
                        p605 = p605 + tc;
                end
                583: begin
                        tc = f582;
                        p607 = p607 - tc;
                        p606 = p606 + tc;
                end
                584: begin
                        tc = f583;
                        p78 = p78 - tc;
                        p603 = p603 + tc;
                        p608 = p608 + tc;
                end
                585: begin
                        tc = f584;
                        p608 = p608 - tc;
                        p78 = p78 + tc;
                end
                586: begin
                        tc = f585;
                        p610 = p610 - tc;
                        p609 = p609 + tc;
                end
                587: begin
                        tc = f586;
                        p611 = p611 - tc;
                        p610 = p610 + tc;
                end
                588: begin
                        tc = f587;
                        p81 = p81 - tc;
                        p604 = p604 + tc;
                        p612 = p612 + tc;
                end
                589: begin
                        tc = f588;
                        p612 = p612 - tc;
                        p81 = p81 + tc;
                end
                590: begin
                        tc = f589;
                        p614 = p614 - tc;
                        p613 = p613 + tc;
                end
                591: begin
                        tc = f590;
                        p615 = p615 - tc;
                        p614 = p614 + tc;
                end
                592: begin
                        tc = f591;
                        p609 = p609 - tc;
                        p613 = p613 - tc;
                        p72 = p72 + tc;
                end
                593: begin
                        tc = f592;
                        p606 = p606 - tc;
                        p611 = p611 + tc;
                        p615 = p615 + tc;
                end
                594: begin
                        tc = f593;
                        p605 = p605 - tc;
                        p82 = p82 + tc;
                end
                595: begin
                        tc = f594;
                        p82 = p82 - tc;
                end
                596: begin
                        tc = f595;
                        p616 = p616 - tc;
                        p607 = p607 + tc;
                end
                597: begin
                        tc = f596;
                        p73 = p73 - tc;
                        p616 = p616 + tc;
                end
                598: begin
                        tc = f597;
                        p623 = p623 - tc;
                        p619 = p619 + tc;
                end
                599: begin
                        tc = f598;
                        p617 = p617 - tc;
                end
                600: begin
                        tc = f599;
                        p621 = p621 - tc;
                        p623 = p623 + tc;
                end
                601: begin
                        tc = f600;
                        p618 = p618 - tc*2;
                        p624 = p624 + tc;
                end
                602: begin
                        tc = f601;
                        p625 = p625 - tc;
                        p622 = p622 + tc;
                end
                603: begin
                        tc = f602;
                        p618 = p618 - tc;
                        p627 = p627 - tc;
                        p626 = p626 + tc;
                end
                604: begin
                        tc = f603;
                        p628 = p628 - tc;
                        p625 = p625 + tc;
                end
                605: begin
                        tc = f604;
                        p617 = p617 - tc;
                        p620 = p620 + tc;
                        p629 = p629 + tc;
                end
                606: begin
                        tc = f605;
                        p617 = p617 - tc;
                        p629 = p629 + tc;
                end
                607: begin
                        tc = f606;
                        p630 = p630 - tc;
                        p628 = p628 + tc;
                end
                608: begin
                        tc = f607;
                        p624 = p624 - tc;
                        p618 = p618 + tc;
                end
                609: begin
                        tc = f608;
                        p631 = p631 - tc;
                        p630 = p630 + tc;
                end
                610: begin
                        tc = f609;
                        p629 = p629 - tc;
                        p617 = p617 + tc*2;
                end
                611: begin
                        tc = f610;
                        p619 = p619 - tc;
                        p626 = p626 - tc;
                        p627 = p627 + tc;
                        p631 = p631 + tc;
                end
                612: begin
                        tc = f611;
                        p619 = p619 - tc;
                        p631 = p631 + tc;
                end
                613: begin
                        tc = f612;
                        p83 = p83 - tc;
                        p617 = p617 + tc;
                        p632 = p632 + tc;
                end
                614: begin
                        tc = f613;
                        p632 = p632 - tc;
                        p83 = p83 + tc;
                end
                615: begin
                        tc = f614;
                        p634 = p634 - tc;
                        p633 = p633 + tc;
                end
                616: begin
                        tc = f615;
                        p635 = p635 - tc;
                        p634 = p634 + tc;
                end
                617: begin
                        tc = f616;
                        p84 = p84 - tc;
                        p618 = p618 + tc;
                        p636 = p636 + tc;
                end
                618: begin
                        tc = f617;
                        p636 = p636 - tc;
                        p84 = p84 + tc;
                end
                619: begin
                        tc = f618;
                        p638 = p638 - tc;
                        p637 = p637 + tc;
                end
                620: begin
                        tc = f619;
                        p639 = p639 - tc;
                        p638 = p638 + tc;
                end
                621: begin
                        tc = f620;
                        p633 = p633 - tc;
                        p637 = p637 - tc;
                        p73 = p73 + tc;
                end
                622: begin
                        tc = f621;
                        p619 = p619 - tc;
                        p635 = p635 + tc;
                        p639 = p639 + tc;
                end
                623: begin
                        tc = f622;
                        p620 = p620 - tc;
                        p85 = p85 + tc;
                end
                624: begin
                        tc = f623;
                        p85 = p85 - tc;
                end
                625: begin
                        tc = f624;
                        p640 = p640 - tc;
                        p621 = p621 + tc;
                end
                626: begin
                        tc = f625;
                        p74 = p74 - tc;
                        p640 = p640 + tc;
                end
                627: begin
                        tc = f626;
                        p642 = p642 - tc;
                        p643 = p643 + tc;
                end
                628: begin
                        tc = f627;
                        p645 = p645 - tc;
                        p644 = p644 + tc;
                end
                629: begin
                        tc = f628;
                        p82 = p82 - tc;
                        p641 = p641 + tc;
                        p646 = p646 + tc;
                end
                630: begin
                        tc = f629;
                        p646 = p646 - tc;
                        p82 = p82 + tc;
                end
                631: begin
                        tc = f630;
                        p648 = p648 - tc;
                        p647 = p647 + tc;
                end
                632: begin
                        tc = f631;
                        p649 = p649 - tc;
                        p648 = p648 + tc;
                end
                633: begin
                        tc = f632;
                        p85 = p85 - tc;
                        p642 = p642 + tc;
                        p650 = p650 + tc;
                end
                634: begin
                        tc = f633;
                        p650 = p650 - tc;
                        p85 = p85 + tc;
                end
                635: begin
                        tc = f634;
                        p652 = p652 - tc;
                        p651 = p651 + tc;
                end
                636: begin
                        tc = f635;
                        p653 = p653 - tc;
                        p652 = p652 + tc;
                end
                637: begin
                        tc = f636;
                        p647 = p647 - tc;
                        p651 = p651 - tc;
                        p74 = p74 + tc;
                end
                638: begin
                        tc = f637;
                        p644 = p644 - tc;
                        p649 = p649 + tc;
                        p653 = p653 + tc;
                end
                639: begin
                        tc = f638;
                        p643 = p643 - tc;
                        p86 = p86 + tc;
                end
                640: begin
                        tc = f639;
                        p86 = p86 - tc;
                end
                641: begin
                        tc = f640;
                        p654 = p654 - tc;
                        p645 = p645 + tc;
                end
                642: begin
                        tc = f641;
                        p75 = p75 - tc;
                        p654 = p654 + tc;
                end
                643: begin
                        tc = f642;
                        p661 = p661 - tc;
                        p657 = p657 + tc;
                end
                644: begin
                        tc = f643;
                        p655 = p655 - tc;
                end
                645: begin
                        tc = f644;
                        p659 = p659 - tc;
                        p661 = p661 + tc;
                end
                646: begin
                        tc = f645;
                        p656 = p656 - tc*2;
                        p662 = p662 + tc;
                end
                647: begin
                        tc = f646;
                        p663 = p663 - tc;
                        p660 = p660 + tc;
                end
                648: begin
                        tc = f647;
                        p656 = p656 - tc;
                        p665 = p665 - tc;
                        p664 = p664 + tc;
                end
                649: begin
                        tc = f648;
                        p666 = p666 - tc;
                        p663 = p663 + tc;
                end
                650: begin
                        tc = f649;
                        p655 = p655 - tc;
                        p658 = p658 + tc;
                        p667 = p667 + tc;
                end
                651: begin
                        tc = f650;
                        p655 = p655 - tc;
                        p667 = p667 + tc;
                end
                652: begin
                        tc = f651;
                        p668 = p668 - tc;
                        p666 = p666 + tc;
                end
                653: begin
                        tc = f652;
                        p662 = p662 - tc;
                        p656 = p656 + tc;
                end
                654: begin
                        tc = f653;
                        p669 = p669 - tc;
                        p668 = p668 + tc;
                end
                655: begin
                        tc = f654;
                        p667 = p667 - tc;
                        p655 = p655 + tc*2;
                end
                656: begin
                        tc = f655;
                        p657 = p657 - tc;
                        p664 = p664 - tc;
                        p665 = p665 + tc;
                        p669 = p669 + tc;
                end
                657: begin
                        tc = f656;
                        p657 = p657 - tc;
                        p669 = p669 + tc;
                end
                658: begin
                        tc = f657;
                        p93 = p93 - tc;
                        p655 = p655 + tc;
                        p670 = p670 + tc;
                end
                659: begin
                        tc = f658;
                        p670 = p670 - tc;
                        p93 = p93 + tc;
                end
                660: begin
                        tc = f659;
                        p672 = p672 - tc;
                        p671 = p671 + tc;
                end
                661: begin
                        tc = f660;
                        p673 = p673 - tc;
                        p672 = p672 + tc;
                end
                662: begin
                        tc = f661;
                        p94 = p94 - tc;
                        p656 = p656 + tc;
                        p674 = p674 + tc;
                end
                663: begin
                        tc = f662;
                        p674 = p674 - tc;
                        p94 = p94 + tc;
                end
                664: begin
                        tc = f663;
                        p676 = p676 - tc;
                        p675 = p675 + tc;
                end
                665: begin
                        tc = f664;
                        p677 = p677 - tc;
                        p676 = p676 + tc;
                end
                666: begin
                        tc = f665;
                        p671 = p671 - tc;
                        p675 = p675 - tc;
                        p87 = p87 + tc;
                end
                667: begin
                        tc = f666;
                        p657 = p657 - tc;
                        p673 = p673 + tc;
                        p677 = p677 + tc;
                end
                668: begin
                        tc = f667;
                        p658 = p658 - tc;
                        p95 = p95 + tc;
                end
                669: begin
                        tc = f668;
                        p95 = p95 - tc;
                end
                670: begin
                        tc = f669;
                        p678 = p678 - tc;
                        p659 = p659 + tc;
                end
                671: begin
                        tc = f670;
                        p88 = p88 - tc;
                        p678 = p678 + tc;
                end
                672: begin
                        tc = f671;
                        p685 = p685 - tc;
                        p681 = p681 + tc;
                end
                673: begin
                        tc = f672;
                        p679 = p679 - tc;
                end
                674: begin
                        tc = f673;
                        p683 = p683 - tc;
                        p685 = p685 + tc;
                end
                675: begin
                        tc = f674;
                        p680 = p680 - tc*2;
                        p686 = p686 + tc;
                end
                676: begin
                        tc = f675;
                        p687 = p687 - tc;
                        p684 = p684 + tc;
                end
                677: begin
                        tc = f676;
                        p680 = p680 - tc;
                        p689 = p689 - tc;
                        p688 = p688 + tc;
                end
                678: begin
                        tc = f677;
                        p690 = p690 - tc;
                        p687 = p687 + tc;
                end
                679: begin
                        tc = f678;
                        p679 = p679 - tc;
                        p682 = p682 + tc;
                        p691 = p691 + tc;
                end
                680: begin
                        tc = f679;
                        p679 = p679 - tc;
                        p691 = p691 + tc;
                end
                681: begin
                        tc = f680;
                        p692 = p692 - tc;
                        p690 = p690 + tc;
                end
                682: begin
                        tc = f681;
                        p686 = p686 - tc;
                        p680 = p680 + tc;
                end
                683: begin
                        tc = f682;
                        p693 = p693 - tc;
                        p692 = p692 + tc;
                end
                684: begin
                        tc = f683;
                        p691 = p691 - tc;
                        p679 = p679 + tc*2;
                end
                685: begin
                        tc = f684;
                        p681 = p681 - tc;
                        p688 = p688 - tc;
                        p689 = p689 + tc;
                        p693 = p693 + tc;
                end
                686: begin
                        tc = f685;
                        p681 = p681 - tc;
                        p693 = p693 + tc;
                end
                687: begin
                        tc = f686;
                        p96 = p96 - tc;
                        p679 = p679 + tc;
                        p694 = p694 + tc;
                end
                688: begin
                        tc = f687;
                        p694 = p694 - tc;
                        p96 = p96 + tc;
                end
                689: begin
                        tc = f688;
                        p696 = p696 - tc;
                        p695 = p695 + tc;
                end
                690: begin
                        tc = f689;
                        p697 = p697 - tc;
                        p696 = p696 + tc;
                end
                691: begin
                        tc = f690;
                        p97 = p97 - tc;
                        p680 = p680 + tc;
                        p698 = p698 + tc;
                end
                692: begin
                        tc = f691;
                        p698 = p698 - tc;
                        p97 = p97 + tc;
                end
                693: begin
                        tc = f692;
                        p700 = p700 - tc;
                        p699 = p699 + tc;
                end
                694: begin
                        tc = f693;
                        p701 = p701 - tc;
                        p700 = p700 + tc;
                end
                695: begin
                        tc = f694;
                        p695 = p695 - tc;
                        p699 = p699 - tc;
                        p88 = p88 + tc;
                end
                696: begin
                        tc = f695;
                        p681 = p681 - tc;
                        p697 = p697 + tc;
                        p701 = p701 + tc;
                end
                697: begin
                        tc = f696;
                        p682 = p682 - tc;
                        p98 = p98 + tc;
                end
                698: begin
                        tc = f697;
                        p98 = p98 - tc;
                end
                699: begin
                        tc = f698;
                        p702 = p702 - tc;
                        p683 = p683 + tc;
                end
                700: begin
                        tc = f699;
                        p89 = p89 - tc;
                        p702 = p702 + tc;
                end
                701: begin
                        tc = f700;
                        p704 = p704 - tc;
                        p705 = p705 + tc;
                end
                702: begin
                        tc = f701;
                        p707 = p707 - tc;
                        p706 = p706 + tc;
                end
                703: begin
                        tc = f702;
                        p95 = p95 - tc;
                        p703 = p703 + tc;
                        p708 = p708 + tc;
                end
                704: begin
                        tc = f703;
                        p708 = p708 - tc;
                        p95 = p95 + tc;
                end
                705: begin
                        tc = f704;
                        p710 = p710 - tc;
                        p709 = p709 + tc;
                end
                706: begin
                        tc = f705;
                        p711 = p711 - tc;
                        p710 = p710 + tc;
                end
                707: begin
                        tc = f706;
                        p98 = p98 - tc;
                        p704 = p704 + tc;
                        p712 = p712 + tc;
                end
                708: begin
                        tc = f707;
                        p712 = p712 - tc;
                        p98 = p98 + tc;
                end
                709: begin
                        tc = f708;
                        p714 = p714 - tc;
                        p713 = p713 + tc;
                end
                710: begin
                        tc = f709;
                        p715 = p715 - tc;
                        p714 = p714 + tc;
                end
                711: begin
                        tc = f710;
                        p709 = p709 - tc;
                        p713 = p713 - tc;
                        p89 = p89 + tc;
                end
                712: begin
                        tc = f711;
                        p706 = p706 - tc;
                        p711 = p711 + tc;
                        p715 = p715 + tc;
                end
                713: begin
                        tc = f712;
                        p705 = p705 - tc;
                        p99 = p99 + tc;
                end
                714: begin
                        tc = f713;
                        p99 = p99 - tc;
                end
                715: begin
                        tc = f714;
                        p716 = p716 - tc;
                        p707 = p707 + tc;
                end
                716: begin
                        tc = f715;
                        p90 = p90 - tc;
                        p716 = p716 + tc;
                end
                717: begin
                        tc = f716;
                        p723 = p723 - tc;
                        p719 = p719 + tc;
                end
                718: begin
                        tc = f717;
                        p717 = p717 - tc;
                end
                719: begin
                        tc = f718;
                        p721 = p721 - tc;
                        p723 = p723 + tc;
                end
                720: begin
                        tc = f719;
                        p718 = p718 - tc*2;
                        p724 = p724 + tc;
                end
                721: begin
                        tc = f720;
                        p725 = p725 - tc;
                        p722 = p722 + tc;
                end
                722: begin
                        tc = f721;
                        p718 = p718 - tc;
                        p727 = p727 - tc;
                        p726 = p726 + tc;
                end
                723: begin
                        tc = f722;
                        p728 = p728 - tc;
                        p725 = p725 + tc;
                end
                724: begin
                        tc = f723;
                        p717 = p717 - tc;
                        p720 = p720 + tc;
                        p729 = p729 + tc;
                end
                725: begin
                        tc = f724;
                        p717 = p717 - tc;
                        p729 = p729 + tc;
                end
                726: begin
                        tc = f725;
                        p730 = p730 - tc;
                        p728 = p728 + tc;
                end
                727: begin
                        tc = f726;
                        p724 = p724 - tc;
                        p718 = p718 + tc;
                end
                728: begin
                        tc = f727;
                        p731 = p731 - tc;
                        p730 = p730 + tc;
                end
                729: begin
                        tc = f728;
                        p729 = p729 - tc;
                        p717 = p717 + tc*2;
                end
                730: begin
                        tc = f729;
                        p719 = p719 - tc;
                        p726 = p726 - tc;
                        p727 = p727 + tc;
                        p731 = p731 + tc;
                end
                731: begin
                        tc = f730;
                        p719 = p719 - tc;
                        p731 = p731 + tc;
                end
                732: begin
                        tc = f731;
                        p100 = p100 - tc;
                        p717 = p717 + tc;
                        p732 = p732 + tc;
                end
                733: begin
                        tc = f732;
                        p732 = p732 - tc;
                        p100 = p100 + tc;
                end
                734: begin
                        tc = f733;
                        p734 = p734 - tc;
                        p733 = p733 + tc;
                end
                735: begin
                        tc = f734;
                        p735 = p735 - tc;
                        p734 = p734 + tc;
                end
                736: begin
                        tc = f735;
                        p101 = p101 - tc;
                        p718 = p718 + tc;
                        p736 = p736 + tc;
                end
                737: begin
                        tc = f736;
                        p736 = p736 - tc;
                        p101 = p101 + tc;
                end
                738: begin
                        tc = f737;
                        p738 = p738 - tc;
                        p737 = p737 + tc;
                end
                739: begin
                        tc = f738;
                        p739 = p739 - tc;
                        p738 = p738 + tc;
                end
                740: begin
                        tc = f739;
                        p733 = p733 - tc;
                        p737 = p737 - tc;
                        p90 = p90 + tc;
                end
                741: begin
                        tc = f740;
                        p719 = p719 - tc;
                        p735 = p735 + tc;
                        p739 = p739 + tc;
                end
                742: begin
                        tc = f741;
                        p720 = p720 - tc;
                        p102 = p102 + tc;
                end
                743: begin
                        tc = f742;
                        p102 = p102 - tc;
                end
                744: begin
                        tc = f743;
                        p740 = p740 - tc;
                        p721 = p721 + tc;
                end
                745: begin
                        tc = f744;
                        p91 = p91 - tc;
                        p740 = p740 + tc;
                end
                746: begin
                        tc = f745;
                        p742 = p742 - tc;
                        p743 = p743 + tc;
                end
                747: begin
                        tc = f746;
                        p745 = p745 - tc;
                        p744 = p744 + tc;
                end
                748: begin
                        tc = f747;
                        p99 = p99 - tc;
                        p741 = p741 + tc;
                        p746 = p746 + tc;
                end
                749: begin
                        tc = f748;
                        p746 = p746 - tc;
                        p99 = p99 + tc;
                end
                750: begin
                        tc = f749;
                        p748 = p748 - tc;
                        p747 = p747 + tc;
                end
                751: begin
                        tc = f750;
                        p749 = p749 - tc;
                        p748 = p748 + tc;
                end
                752: begin
                        tc = f751;
                        p102 = p102 - tc;
                        p742 = p742 + tc;
                        p750 = p750 + tc;
                end
                753: begin
                        tc = f752;
                        p750 = p750 - tc;
                        p102 = p102 + tc;
                end
                754: begin
                        tc = f753;
                        p752 = p752 - tc;
                        p751 = p751 + tc;
                end
                755: begin
                        tc = f754;
                        p753 = p753 - tc;
                        p752 = p752 + tc;
                end
                756: begin
                        tc = f755;
                        p747 = p747 - tc;
                        p751 = p751 - tc;
                        p91 = p91 + tc;
                end
                757: begin
                        tc = f756;
                        p744 = p744 - tc;
                        p749 = p749 + tc;
                        p753 = p753 + tc;
                end
                758: begin
                        tc = f757;
                        p743 = p743 - tc;
                        p103 = p103 + tc;
                end
                759: begin
                        tc = f758;
                        p103 = p103 - tc;
                end
                760: begin
                        tc = f759;
                        p754 = p754 - tc;
                        p745 = p745 + tc;
                end
                761: begin
                        tc = f760;
                        p92 = p92 - tc;
                        p754 = p754 + tc;
                end
                762: begin
                        tc = f761;
                        p761 = p761 - tc;
                        p757 = p757 + tc;
                end
                763: begin
                        tc = f762;
                        p755 = p755 - tc;
                end
                764: begin
                        tc = f763;
                        p759 = p759 - tc;
                        p761 = p761 + tc;
                end
                765: begin
                        tc = f764;
                        p756 = p756 - tc*2;
                        p762 = p762 + tc;
                end
                766: begin
                        tc = f765;
                        p763 = p763 - tc;
                        p760 = p760 + tc;
                end
                767: begin
                        tc = f766;
                        p756 = p756 - tc;
                        p765 = p765 - tc;
                        p764 = p764 + tc;
                end
                768: begin
                        tc = f767;
                        p766 = p766 - tc;
                        p763 = p763 + tc;
                end
                769: begin
                        tc = f768;
                        p755 = p755 - tc;
                        p758 = p758 + tc;
                        p767 = p767 + tc;
                end
                770: begin
                        tc = f769;
                        p755 = p755 - tc;
                        p767 = p767 + tc;
                end
                771: begin
                        tc = f770;
                        p768 = p768 - tc;
                        p766 = p766 + tc;
                end
                772: begin
                        tc = f771;
                        p762 = p762 - tc;
                        p756 = p756 + tc;
                end
                773: begin
                        tc = f772;
                        p769 = p769 - tc;
                        p768 = p768 + tc;
                end
                774: begin
                        tc = f773;
                        p767 = p767 - tc;
                        p755 = p755 + tc*2;
                end
                775: begin
                        tc = f774;
                        p757 = p757 - tc;
                        p764 = p764 - tc;
                        p765 = p765 + tc;
                        p769 = p769 + tc;
                end
                776: begin
                        tc = f775;
                        p757 = p757 - tc;
                        p769 = p769 + tc;
                end
                777: begin
                        tc = f776;
                        p110 = p110 - tc;
                        p755 = p755 + tc;
                        p770 = p770 + tc;
                end
                778: begin
                        tc = f777;
                        p770 = p770 - tc;
                        p110 = p110 + tc;
                end
                779: begin
                        tc = f778;
                        p772 = p772 - tc;
                        p771 = p771 + tc;
                end
                780: begin
                        tc = f779;
                        p773 = p773 - tc;
                        p772 = p772 + tc;
                end
                781: begin
                        tc = f780;
                        p111 = p111 - tc;
                        p756 = p756 + tc;
                        p774 = p774 + tc;
                end
                782: begin
                        tc = f781;
                        p774 = p774 - tc;
                        p111 = p111 + tc;
                end
                783: begin
                        tc = f782;
                        p776 = p776 - tc;
                        p775 = p775 + tc;
                end
                784: begin
                        tc = f783;
                        p777 = p777 - tc;
                        p776 = p776 + tc;
                end
                785: begin
                        tc = f784;
                        p771 = p771 - tc;
                        p775 = p775 - tc;
                        p104 = p104 + tc;
                end
                786: begin
                        tc = f785;
                        p757 = p757 - tc;
                        p773 = p773 + tc;
                        p777 = p777 + tc;
                end
                787: begin
                        tc = f786;
                        p758 = p758 - tc;
                        p112 = p112 + tc;
                end
                788: begin
                        tc = f787;
                        p112 = p112 - tc;
                end
                789: begin
                        tc = f788;
                        p778 = p778 - tc;
                        p759 = p759 + tc;
                end
                790: begin
                        tc = f789;
                        p105 = p105 - tc;
                        p778 = p778 + tc;
                end
                791: begin
                        tc = f790;
                        p785 = p785 - tc;
                        p781 = p781 + tc;
                end
                792: begin
                        tc = f791;
                        p779 = p779 - tc;
                end
                793: begin
                        tc = f792;
                        p783 = p783 - tc;
                        p785 = p785 + tc;
                end
                794: begin
                        tc = f793;
                        p780 = p780 - tc*2;
                        p786 = p786 + tc;
                end
                795: begin
                        tc = f794;
                        p787 = p787 - tc;
                        p784 = p784 + tc;
                end
                796: begin
                        tc = f795;
                        p780 = p780 - tc;
                        p789 = p789 - tc;
                        p788 = p788 + tc;
                end
                797: begin
                        tc = f796;
                        p790 = p790 - tc;
                        p787 = p787 + tc;
                end
                798: begin
                        tc = f797;
                        p779 = p779 - tc;
                        p782 = p782 + tc;
                        p791 = p791 + tc;
                end
                799: begin
                        tc = f798;
                        p779 = p779 - tc;
                        p791 = p791 + tc;
                end
                800: begin
                        tc = f799;
                        p792 = p792 - tc;
                        p790 = p790 + tc;
                end
                801: begin
                        tc = f800;
                        p786 = p786 - tc;
                        p780 = p780 + tc;
                end
                802: begin
                        tc = f801;
                        p793 = p793 - tc;
                        p792 = p792 + tc;
                end
                803: begin
                        tc = f802;
                        p791 = p791 - tc;
                        p779 = p779 + tc*2;
                end
                804: begin
                        tc = f803;
                        p781 = p781 - tc;
                        p788 = p788 - tc;
                        p789 = p789 + tc;
                        p793 = p793 + tc;
                end
                805: begin
                        tc = f804;
                        p781 = p781 - tc;
                        p793 = p793 + tc;
                end
                806: begin
                        tc = f805;
                        p113 = p113 - tc;
                        p779 = p779 + tc;
                        p794 = p794 + tc;
                end
                807: begin
                        tc = f806;
                        p794 = p794 - tc;
                        p113 = p113 + tc;
                end
                808: begin
                        tc = f807;
                        p796 = p796 - tc;
                        p795 = p795 + tc;
                end
                809: begin
                        tc = f808;
                        p797 = p797 - tc;
                        p796 = p796 + tc;
                end
                810: begin
                        tc = f809;
                        p114 = p114 - tc;
                        p780 = p780 + tc;
                        p798 = p798 + tc;
                end
                811: begin
                        tc = f810;
                        p798 = p798 - tc;
                        p114 = p114 + tc;
                end
                812: begin
                        tc = f811;
                        p800 = p800 - tc;
                        p799 = p799 + tc;
                end
                813: begin
                        tc = f812;
                        p801 = p801 - tc;
                        p800 = p800 + tc;
                end
                814: begin
                        tc = f813;
                        p795 = p795 - tc;
                        p799 = p799 - tc;
                        p105 = p105 + tc;
                end
                815: begin
                        tc = f814;
                        p781 = p781 - tc;
                        p797 = p797 + tc;
                        p801 = p801 + tc;
                end
                816: begin
                        tc = f815;
                        p782 = p782 - tc;
                        p115 = p115 + tc;
                end
                817: begin
                        tc = f816;
                        p115 = p115 - tc;
                end
                818: begin
                        tc = f817;
                        p802 = p802 - tc;
                        p783 = p783 + tc;
                end
                819: begin
                        tc = f818;
                        p106 = p106 - tc;
                        p802 = p802 + tc;
                end
                820: begin
                        tc = f819;
                        p804 = p804 - tc;
                        p805 = p805 + tc;
                end
                821: begin
                        tc = f820;
                        p807 = p807 - tc;
                        p806 = p806 + tc;
                end
                822: begin
                        tc = f821;
                        p112 = p112 - tc;
                        p803 = p803 + tc;
                        p808 = p808 + tc;
                end
                823: begin
                        tc = f822;
                        p808 = p808 - tc;
                        p112 = p112 + tc;
                end
                824: begin
                        tc = f823;
                        p810 = p810 - tc;
                        p809 = p809 + tc;
                end
                825: begin
                        tc = f824;
                        p811 = p811 - tc;
                        p810 = p810 + tc;
                end
                826: begin
                        tc = f825;
                        p115 = p115 - tc;
                        p804 = p804 + tc;
                        p812 = p812 + tc;
                end
                827: begin
                        tc = f826;
                        p812 = p812 - tc;
                        p115 = p115 + tc;
                end
                828: begin
                        tc = f827;
                        p814 = p814 - tc;
                        p813 = p813 + tc;
                end
                829: begin
                        tc = f828;
                        p815 = p815 - tc;
                        p814 = p814 + tc;
                end
                830: begin
                        tc = f829;
                        p809 = p809 - tc;
                        p813 = p813 - tc;
                        p106 = p106 + tc;
                end
                831: begin
                        tc = f830;
                        p806 = p806 - tc;
                        p811 = p811 + tc;
                        p815 = p815 + tc;
                end
                832: begin
                        tc = f831;
                        p805 = p805 - tc;
                        p116 = p116 + tc;
                end
                833: begin
                        tc = f832;
                        p116 = p116 - tc;
                end
                834: begin
                        tc = f833;
                        p816 = p816 - tc;
                        p807 = p807 + tc;
                end
                835: begin
                        tc = f834;
                        p107 = p107 - tc;
                        p816 = p816 + tc;
                end
                836: begin
                        tc = f835;
                        p823 = p823 - tc;
                        p819 = p819 + tc;
                end
                837: begin
                        tc = f836;
                        p817 = p817 - tc;
                end
                838: begin
                        tc = f837;
                        p821 = p821 - tc;
                        p823 = p823 + tc;
                end
                839: begin
                        tc = f838;
                        p818 = p818 - tc*2;
                        p824 = p824 + tc;
                end
                840: begin
                        tc = f839;
                        p825 = p825 - tc;
                        p822 = p822 + tc;
                end
                841: begin
                        tc = f840;
                        p818 = p818 - tc;
                        p827 = p827 - tc;
                        p826 = p826 + tc;
                end
                842: begin
                        tc = f841;
                        p828 = p828 - tc;
                        p825 = p825 + tc;
                end
                843: begin
                        tc = f842;
                        p817 = p817 - tc;
                        p820 = p820 + tc;
                        p829 = p829 + tc;
                end
                844: begin
                        tc = f843;
                        p817 = p817 - tc;
                        p829 = p829 + tc;
                end
                845: begin
                        tc = f844;
                        p830 = p830 - tc;
                        p828 = p828 + tc;
                end
                846: begin
                        tc = f845;
                        p824 = p824 - tc;
                        p818 = p818 + tc;
                end
                847: begin
                        tc = f846;
                        p831 = p831 - tc;
                        p830 = p830 + tc;
                end
                848: begin
                        tc = f847;
                        p829 = p829 - tc;
                        p817 = p817 + tc*2;
                end
                849: begin
                        tc = f848;
                        p819 = p819 - tc;
                        p826 = p826 - tc;
                        p827 = p827 + tc;
                        p831 = p831 + tc;
                end
                850: begin
                        tc = f849;
                        p819 = p819 - tc;
                        p831 = p831 + tc;
                end
                851: begin
                        tc = f850;
                        p117 = p117 - tc;
                        p817 = p817 + tc;
                        p832 = p832 + tc;
                end
                852: begin
                        tc = f851;
                        p832 = p832 - tc;
                        p117 = p117 + tc;
                end
                853: begin
                        tc = f852;
                        p834 = p834 - tc;
                        p833 = p833 + tc;
                end
                854: begin
                        tc = f853;
                        p835 = p835 - tc;
                        p834 = p834 + tc;
                end
                855: begin
                        tc = f854;
                        p118 = p118 - tc;
                        p818 = p818 + tc;
                        p836 = p836 + tc;
                end
                856: begin
                        tc = f855;
                        p836 = p836 - tc;
                        p118 = p118 + tc;
                end
                857: begin
                        tc = f856;
                        p838 = p838 - tc;
                        p837 = p837 + tc;
                end
                858: begin
                        tc = f857;
                        p839 = p839 - tc;
                        p838 = p838 + tc;
                end
                859: begin
                        tc = f858;
                        p833 = p833 - tc;
                        p837 = p837 - tc;
                        p107 = p107 + tc;
                end
                860: begin
                        tc = f859;
                        p819 = p819 - tc;
                        p835 = p835 + tc;
                        p839 = p839 + tc;
                end
                861: begin
                        tc = f860;
                        p820 = p820 - tc;
                        p119 = p119 + tc;
                end
                862: begin
                        tc = f861;
                        p119 = p119 - tc;
                end
                863: begin
                        tc = f862;
                        p840 = p840 - tc;
                        p821 = p821 + tc;
                end
                864: begin
                        tc = f863;
                        p108 = p108 - tc;
                        p840 = p840 + tc;
                end
                865: begin
                        tc = f864;
                        p842 = p842 - tc;
                        p843 = p843 + tc;
                end
                866: begin
                        tc = f865;
                        p845 = p845 - tc;
                        p844 = p844 + tc;
                end
                867: begin
                        tc = f866;
                        p116 = p116 - tc;
                        p841 = p841 + tc;
                        p846 = p846 + tc;
                end
                868: begin
                        tc = f867;
                        p846 = p846 - tc;
                        p116 = p116 + tc;
                end
                869: begin
                        tc = f868;
                        p848 = p848 - tc;
                        p847 = p847 + tc;
                end
                870: begin
                        tc = f869;
                        p849 = p849 - tc;
                        p848 = p848 + tc;
                end
                871: begin
                        tc = f870;
                        p119 = p119 - tc;
                        p842 = p842 + tc;
                        p850 = p850 + tc;
                end
                872: begin
                        tc = f871;
                        p850 = p850 - tc;
                        p119 = p119 + tc;
                end
                873: begin
                        tc = f872;
                        p852 = p852 - tc;
                        p851 = p851 + tc;
                end
                874: begin
                        tc = f873;
                        p853 = p853 - tc;
                        p852 = p852 + tc;
                end
                875: begin
                        tc = f874;
                        p847 = p847 - tc;
                        p851 = p851 - tc;
                        p108 = p108 + tc;
                end
                876: begin
                        tc = f875;
                        p844 = p844 - tc;
                        p849 = p849 + tc;
                        p853 = p853 + tc;
                end
                877: begin
                        tc = f876;
                        p843 = p843 - tc;
                        p120 = p120 + tc;
                end
                878: begin
                        tc = f877;
                        p120 = p120 - tc;
                end
                879: begin
                        tc = f878;
                        p854 = p854 - tc;
                        p845 = p845 + tc;
                end
                880: begin
                        tc = f879;
                        p109 = p109 - tc;
                        p854 = p854 + tc;
                end
                881: begin
                        tc = f880;
                        p861 = p861 - tc;
                        p857 = p857 + tc;
                end
                882: begin
                        tc = f881;
                        p855 = p855 - tc;
                end
                883: begin
                        tc = f882;
                        p859 = p859 - tc;
                        p861 = p861 + tc;
                end
                884: begin
                        tc = f883;
                        p856 = p856 - tc*2;
                        p862 = p862 + tc;
                end
                885: begin
                        tc = f884;
                        p863 = p863 - tc;
                        p860 = p860 + tc;
                end
                886: begin
                        tc = f885;
                        p856 = p856 - tc;
                        p865 = p865 - tc;
                        p864 = p864 + tc;
                end
                887: begin
                        tc = f886;
                        p866 = p866 - tc;
                        p863 = p863 + tc;
                end
                888: begin
                        tc = f887;
                        p855 = p855 - tc;
                        p858 = p858 + tc;
                        p867 = p867 + tc;
                end
                889: begin
                        tc = f888;
                        p855 = p855 - tc;
                        p867 = p867 + tc;
                end
                890: begin
                        tc = f889;
                        p868 = p868 - tc;
                        p866 = p866 + tc;
                end
                891: begin
                        tc = f890;
                        p862 = p862 - tc;
                        p856 = p856 + tc;
                end
                892: begin
                        tc = f891;
                        p869 = p869 - tc;
                        p868 = p868 + tc;
                end
                893: begin
                        tc = f892;
                        p867 = p867 - tc;
                        p855 = p855 + tc*2;
                end
                894: begin
                        tc = f893;
                        p857 = p857 - tc;
                        p864 = p864 - tc;
                        p865 = p865 + tc;
                        p869 = p869 + tc;
                end
                895: begin
                        tc = f894;
                        p857 = p857 - tc;
                        p869 = p869 + tc;
                end
                896: begin
                        tc = f895;
                        p127 = p127 - tc;
                        p855 = p855 + tc;
                        p870 = p870 + tc;
                end
                897: begin
                        tc = f896;
                        p870 = p870 - tc;
                        p127 = p127 + tc;
                end
                898: begin
                        tc = f897;
                        p872 = p872 - tc;
                        p871 = p871 + tc;
                end
                899: begin
                        tc = f898;
                        p873 = p873 - tc;
                        p872 = p872 + tc;
                end
                900: begin
                        tc = f899;
                        p128 = p128 - tc;
                        p856 = p856 + tc;
                        p874 = p874 + tc;
                end
                901: begin
                        tc = f900;
                        p874 = p874 - tc;
                        p128 = p128 + tc;
                end
                902: begin
                        tc = f901;
                        p876 = p876 - tc;
                        p875 = p875 + tc;
                end
                903: begin
                        tc = f902;
                        p877 = p877 - tc;
                        p876 = p876 + tc;
                end
                904: begin
                        tc = f903;
                        p871 = p871 - tc;
                        p875 = p875 - tc;
                        p121 = p121 + tc;
                end
                905: begin
                        tc = f904;
                        p857 = p857 - tc;
                        p873 = p873 + tc;
                        p877 = p877 + tc;
                end
                906: begin
                        tc = f905;
                        p858 = p858 - tc;
                        p129 = p129 + tc;
                end
                907: begin
                        tc = f906;
                        p129 = p129 - tc;
                end
                908: begin
                        tc = f907;
                        p878 = p878 - tc;
                        p859 = p859 + tc;
                end
                909: begin
                        tc = f908;
                        p122 = p122 - tc;
                        p878 = p878 + tc;
                end
                910: begin
                        tc = f909;
                        p885 = p885 - tc;
                        p881 = p881 + tc;
                end
                911: begin
                        tc = f910;
                        p879 = p879 - tc;
                end
                912: begin
                        tc = f911;
                        p883 = p883 - tc;
                        p885 = p885 + tc;
                end
                913: begin
                        tc = f912;
                        p880 = p880 - tc*2;
                        p886 = p886 + tc;
                end
                914: begin
                        tc = f913;
                        p887 = p887 - tc;
                        p884 = p884 + tc;
                end
                915: begin
                        tc = f914;
                        p880 = p880 - tc;
                        p889 = p889 - tc;
                        p888 = p888 + tc;
                end
                916: begin
                        tc = f915;
                        p890 = p890 - tc;
                        p887 = p887 + tc;
                end
                917: begin
                        tc = f916;
                        p879 = p879 - tc;
                        p882 = p882 + tc;
                        p891 = p891 + tc;
                end
                918: begin
                        tc = f917;
                        p879 = p879 - tc;
                        p891 = p891 + tc;
                end
                919: begin
                        tc = f918;
                        p892 = p892 - tc;
                        p890 = p890 + tc;
                end
                920: begin
                        tc = f919;
                        p886 = p886 - tc;
                        p880 = p880 + tc;
                end
                921: begin
                        tc = f920;
                        p893 = p893 - tc;
                        p892 = p892 + tc;
                end
                922: begin
                        tc = f921;
                        p891 = p891 - tc;
                        p879 = p879 + tc*2;
                end
                923: begin
                        tc = f922;
                        p881 = p881 - tc;
                        p888 = p888 - tc;
                        p889 = p889 + tc;
                        p893 = p893 + tc;
                end
                924: begin
                        tc = f923;
                        p881 = p881 - tc;
                        p893 = p893 + tc;
                end
                925: begin
                        tc = f924;
                        p130 = p130 - tc;
                        p879 = p879 + tc;
                        p894 = p894 + tc;
                end
                926: begin
                        tc = f925;
                        p894 = p894 - tc;
                        p130 = p130 + tc;
                end
                927: begin
                        tc = f926;
                        p896 = p896 - tc;
                        p895 = p895 + tc;
                end
                928: begin
                        tc = f927;
                        p897 = p897 - tc;
                        p896 = p896 + tc;
                end
                929: begin
                        tc = f928;
                        p131 = p131 - tc;
                        p880 = p880 + tc;
                        p898 = p898 + tc;
                end
                930: begin
                        tc = f929;
                        p898 = p898 - tc;
                        p131 = p131 + tc;
                end
                931: begin
                        tc = f930;
                        p900 = p900 - tc;
                        p899 = p899 + tc;
                end
                932: begin
                        tc = f931;
                        p901 = p901 - tc;
                        p900 = p900 + tc;
                end
                933: begin
                        tc = f932;
                        p895 = p895 - tc;
                        p899 = p899 - tc;
                        p122 = p122 + tc;
                end
                934: begin
                        tc = f933;
                        p881 = p881 - tc;
                        p897 = p897 + tc;
                        p901 = p901 + tc;
                end
                935: begin
                        tc = f934;
                        p882 = p882 - tc;
                        p132 = p132 + tc;
                end
                936: begin
                        tc = f935;
                        p132 = p132 - tc;
                end
                937: begin
                        tc = f936;
                        p902 = p902 - tc;
                        p883 = p883 + tc;
                end
                938: begin
                        tc = f937;
                        p123 = p123 - tc;
                        p902 = p902 + tc;
                end
                939: begin
                        tc = f938;
                        p904 = p904 - tc;
                        p905 = p905 + tc;
                end
                940: begin
                        tc = f939;
                        p907 = p907 - tc;
                        p906 = p906 + tc;
                end
                941: begin
                        tc = f940;
                        p129 = p129 - tc;
                        p903 = p903 + tc;
                        p908 = p908 + tc;
                end
                942: begin
                        tc = f941;
                        p908 = p908 - tc;
                        p129 = p129 + tc;
                end
                943: begin
                        tc = f942;
                        p910 = p910 - tc;
                        p909 = p909 + tc;
                end
                944: begin
                        tc = f943;
                        p911 = p911 - tc;
                        p910 = p910 + tc;
                end
                945: begin
                        tc = f944;
                        p132 = p132 - tc;
                        p904 = p904 + tc;
                        p912 = p912 + tc;
                end
                946: begin
                        tc = f945;
                        p912 = p912 - tc;
                        p132 = p132 + tc;
                end
                947: begin
                        tc = f946;
                        p914 = p914 - tc;
                        p913 = p913 + tc;
                end
                948: begin
                        tc = f947;
                        p915 = p915 - tc;
                        p914 = p914 + tc;
                end
                949: begin
                        tc = f948;
                        p909 = p909 - tc;
                        p913 = p913 - tc;
                        p123 = p123 + tc;
                end
                950: begin
                        tc = f949;
                        p906 = p906 - tc;
                        p911 = p911 + tc;
                        p915 = p915 + tc;
                end
                951: begin
                        tc = f950;
                        p905 = p905 - tc;
                        p133 = p133 + tc;
                end
                952: begin
                        tc = f951;
                        p133 = p133 - tc;
                end
                953: begin
                        tc = f952;
                        p916 = p916 - tc;
                        p907 = p907 + tc;
                end
                954: begin
                        tc = f953;
                        p124 = p124 - tc;
                        p916 = p916 + tc;
                end
                955: begin
                        tc = f954;
                        p923 = p923 - tc;
                        p919 = p919 + tc;
                end
                956: begin
                        tc = f955;
                        p917 = p917 - tc;
                end
                957: begin
                        tc = f956;
                        p921 = p921 - tc;
                        p923 = p923 + tc;
                end
                958: begin
                        tc = f957;
                        p918 = p918 - tc*2;
                        p924 = p924 + tc;
                end
                959: begin
                        tc = f958;
                        p925 = p925 - tc;
                        p922 = p922 + tc;
                end
                960: begin
                        tc = f959;
                        p918 = p918 - tc;
                        p927 = p927 - tc;
                        p926 = p926 + tc;
                end
                961: begin
                        tc = f960;
                        p928 = p928 - tc;
                        p925 = p925 + tc;
                end
                962: begin
                        tc = f961;
                        p917 = p917 - tc;
                        p920 = p920 + tc;
                        p929 = p929 + tc;
                end
                963: begin
                        tc = f962;
                        p917 = p917 - tc;
                        p929 = p929 + tc;
                end
                964: begin
                        tc = f963;
                        p930 = p930 - tc;
                        p928 = p928 + tc;
                end
                965: begin
                        tc = f964;
                        p924 = p924 - tc;
                        p918 = p918 + tc;
                end
                966: begin
                        tc = f965;
                        p931 = p931 - tc;
                        p930 = p930 + tc;
                end
                967: begin
                        tc = f966;
                        p929 = p929 - tc;
                        p917 = p917 + tc*2;
                end
                968: begin
                        tc = f967;
                        p919 = p919 - tc;
                        p926 = p926 - tc;
                        p927 = p927 + tc;
                        p931 = p931 + tc;
                end
                969: begin
                        tc = f968;
                        p919 = p919 - tc;
                        p931 = p931 + tc;
                end
                970: begin
                        tc = f969;
                        p134 = p134 - tc;
                        p917 = p917 + tc;
                        p932 = p932 + tc;
                end
                971: begin
                        tc = f970;
                        p932 = p932 - tc;
                        p134 = p134 + tc;
                end
                972: begin
                        tc = f971;
                        p934 = p934 - tc;
                        p933 = p933 + tc;
                end
                973: begin
                        tc = f972;
                        p935 = p935 - tc;
                        p934 = p934 + tc;
                end
                974: begin
                        tc = f973;
                        p135 = p135 - tc;
                        p918 = p918 + tc;
                        p936 = p936 + tc;
                end
                975: begin
                        tc = f974;
                        p936 = p936 - tc;
                        p135 = p135 + tc;
                end
                976: begin
                        tc = f975;
                        p938 = p938 - tc;
                        p937 = p937 + tc;
                end
                977: begin
                        tc = f976;
                        p939 = p939 - tc;
                        p938 = p938 + tc;
                end
                978: begin
                        tc = f977;
                        p933 = p933 - tc;
                        p937 = p937 - tc;
                        p124 = p124 + tc;
                end
                979: begin
                        tc = f978;
                        p919 = p919 - tc;
                        p935 = p935 + tc;
                        p939 = p939 + tc;
                end
                980: begin
                        tc = f979;
                        p920 = p920 - tc;
                        p136 = p136 + tc;
                end
                981: begin
                        tc = f980;
                        p136 = p136 - tc;
                end
                982: begin
                        tc = f981;
                        p940 = p940 - tc;
                        p921 = p921 + tc;
                end
                983: begin
                        tc = f982;
                        p125 = p125 - tc;
                        p940 = p940 + tc;
                end
                984: begin
                        tc = f983;
                        p942 = p942 - tc;
                        p943 = p943 + tc;
                end
                985: begin
                        tc = f984;
                        p945 = p945 - tc;
                        p944 = p944 + tc;
                end
                986: begin
                        tc = f985;
                        p133 = p133 - tc;
                        p941 = p941 + tc;
                        p946 = p946 + tc;
                end
                987: begin
                        tc = f986;
                        p946 = p946 - tc;
                        p133 = p133 + tc;
                end
                988: begin
                        tc = f987;
                        p948 = p948 - tc;
                        p947 = p947 + tc;
                end
                989: begin
                        tc = f988;
                        p949 = p949 - tc;
                        p948 = p948 + tc;
                end
                990: begin
                        tc = f989;
                        p136 = p136 - tc;
                        p942 = p942 + tc;
                        p950 = p950 + tc;
                end
                991: begin
                        tc = f990;
                        p950 = p950 - tc;
                        p136 = p136 + tc;
                end
                992: begin
                        tc = f991;
                        p952 = p952 - tc;
                        p951 = p951 + tc;
                end
                993: begin
                        tc = f992;
                        p953 = p953 - tc;
                        p952 = p952 + tc;
                end
                994: begin
                        tc = f993;
                        p947 = p947 - tc;
                        p951 = p951 - tc;
                        p125 = p125 + tc;
                end
                995: begin
                        tc = f994;
                        p944 = p944 - tc;
                        p949 = p949 + tc;
                        p953 = p953 + tc;
                end
                996: begin
                        tc = f995;
                        p943 = p943 - tc;
                        p137 = p137 + tc;
                end
                997: begin
                        tc = f996;
                        p137 = p137 - tc;
                end
                998: begin
                        tc = f997;
                        p954 = p954 - tc;
                        p945 = p945 + tc;
                end
                999: begin
                        tc = f998;
                        p126 = p126 - tc;
                        p954 = p954 + tc;
                end
                1000: begin
                        tc = f999;
                        p961 = p961 - tc;
                        p957 = p957 + tc;
                end
                1001: begin
                        tc = f1000;
                        p955 = p955 - tc;
                end
                1002: begin
                        tc = f1001;
                        p959 = p959 - tc;
                        p961 = p961 + tc;
                end
                1003: begin
                        tc = f1002;
                        p956 = p956 - tc*2;
                        p962 = p962 + tc;
                end
                1004: begin
                        tc = f1003;
                        p963 = p963 - tc;
                        p960 = p960 + tc;
                end
                1005: begin
                        tc = f1004;
                        p956 = p956 - tc;
                        p965 = p965 - tc;
                        p964 = p964 + tc;
                end
                1006: begin
                        tc = f1005;
                        p966 = p966 - tc;
                        p963 = p963 + tc;
                end
                1007: begin
                        tc = f1006;
                        p955 = p955 - tc;
                        p958 = p958 + tc;
                        p967 = p967 + tc;
                end
                1008: begin
                        tc = f1007;
                        p955 = p955 - tc;
                        p967 = p967 + tc;
                end
                1009: begin
                        tc = f1008;
                        p968 = p968 - tc;
                        p966 = p966 + tc;
                end
                1010: begin
                        tc = f1009;
                        p962 = p962 - tc;
                        p956 = p956 + tc;
                end
                1011: begin
                        tc = f1010;
                        p969 = p969 - tc;
                        p968 = p968 + tc;
                end
                1012: begin
                        tc = f1011;
                        p967 = p967 - tc;
                        p955 = p955 + tc*2;
                end
                1013: begin
                        tc = f1012;
                        p957 = p957 - tc;
                        p964 = p964 - tc;
                        p965 = p965 + tc;
                        p969 = p969 + tc;
                end
                1014: begin
                        tc = f1013;
                        p957 = p957 - tc;
                        p969 = p969 + tc;
                end
                1015: begin
                        tc = f1014;
                        p144 = p144 - tc;
                        p955 = p955 + tc;
                        p970 = p970 + tc;
                end
                1016: begin
                        tc = f1015;
                        p970 = p970 - tc;
                        p144 = p144 + tc;
                end
                1017: begin
                        tc = f1016;
                        p972 = p972 - tc;
                        p971 = p971 + tc;
                end
                1018: begin
                        tc = f1017;
                        p973 = p973 - tc;
                        p972 = p972 + tc;
                end
                1019: begin
                        tc = f1018;
                        p145 = p145 - tc;
                        p956 = p956 + tc;
                        p974 = p974 + tc;
                end
                1020: begin
                        tc = f1019;
                        p974 = p974 - tc;
                        p145 = p145 + tc;
                end
                1021: begin
                        tc = f1020;
                        p976 = p976 - tc;
                        p975 = p975 + tc;
                end
                1022: begin
                        tc = f1021;
                        p977 = p977 - tc;
                        p976 = p976 + tc;
                end
                1023: begin
                        tc = f1022;
                        p971 = p971 - tc;
                        p975 = p975 - tc;
                        p138 = p138 + tc;
                end
                1024: begin
                        tc = f1023;
                        p957 = p957 - tc;
                        p973 = p973 + tc;
                        p977 = p977 + tc;
                end
                1025: begin
                        tc = f1024;
                        p958 = p958 - tc;
                        p146 = p146 + tc;
                end
                1026: begin
                        tc = f1025;
                        p146 = p146 - tc;
                end
                1027: begin
                        tc = f1026;
                        p978 = p978 - tc;
                        p959 = p959 + tc;
                end
                1028: begin
                        tc = f1027;
                        p139 = p139 - tc;
                        p978 = p978 + tc;
                end
                1029: begin
                        tc = f1028;
                        p985 = p985 - tc;
                        p981 = p981 + tc;
                end
                1030: begin
                        tc = f1029;
                        p979 = p979 - tc;
                end
                1031: begin
                        tc = f1030;
                        p983 = p983 - tc;
                        p985 = p985 + tc;
                end
                1032: begin
                        tc = f1031;
                        p980 = p980 - tc*2;
                        p986 = p986 + tc;
                end
                1033: begin
                        tc = f1032;
                        p987 = p987 - tc;
                        p984 = p984 + tc;
                end
                1034: begin
                        tc = f1033;
                        p980 = p980 - tc;
                        p989 = p989 - tc;
                        p988 = p988 + tc;
                end
                1035: begin
                        tc = f1034;
                        p990 = p990 - tc;
                        p987 = p987 + tc;
                end
                1036: begin
                        tc = f1035;
                        p979 = p979 - tc;
                        p982 = p982 + tc;
                        p991 = p991 + tc;
                end
                1037: begin
                        tc = f1036;
                        p979 = p979 - tc;
                        p991 = p991 + tc;
                end
                1038: begin
                        tc = f1037;
                        p992 = p992 - tc;
                        p990 = p990 + tc;
                end
                1039: begin
                        tc = f1038;
                        p986 = p986 - tc;
                        p980 = p980 + tc;
                end
                1040: begin
                        tc = f1039;
                        p993 = p993 - tc;
                        p992 = p992 + tc;
                end
                1041: begin
                        tc = f1040;
                        p991 = p991 - tc;
                        p979 = p979 + tc*2;
                end
                1042: begin
                        tc = f1041;
                        p981 = p981 - tc;
                        p988 = p988 - tc;
                        p989 = p989 + tc;
                        p993 = p993 + tc;
                end
                1043: begin
                        tc = f1042;
                        p981 = p981 - tc;
                        p993 = p993 + tc;
                end
                1044: begin
                        tc = f1043;
                        p147 = p147 - tc;
                        p979 = p979 + tc;
                        p994 = p994 + tc;
                end
                1045: begin
                        tc = f1044;
                        p994 = p994 - tc;
                        p147 = p147 + tc;
                end
                1046: begin
                        tc = f1045;
                        p996 = p996 - tc;
                        p995 = p995 + tc;
                end
                1047: begin
                        tc = f1046;
                        p997 = p997 - tc;
                        p996 = p996 + tc;
                end
                1048: begin
                        tc = f1047;
                        p148 = p148 - tc;
                        p980 = p980 + tc;
                        p998 = p998 + tc;
                end
                1049: begin
                        tc = f1048;
                        p998 = p998 - tc;
                        p148 = p148 + tc;
                end
                1050: begin
                        tc = f1049;
                        p1000 = p1000 - tc;
                        p999 = p999 + tc;
                end
                1051: begin
                        tc = f1050;
                        p1001 = p1001 - tc;
                        p1000 = p1000 + tc;
                end
                1052: begin
                        tc = f1051;
                        p995 = p995 - tc;
                        p999 = p999 - tc;
                        p139 = p139 + tc;
                end
                1053: begin
                        tc = f1052;
                        p981 = p981 - tc;
                        p997 = p997 + tc;
                        p1001 = p1001 + tc;
                end
                1054: begin
                        tc = f1053;
                        p982 = p982 - tc;
                        p149 = p149 + tc;
                end
                1055: begin
                        tc = f1054;
                        p149 = p149 - tc;
                end
                1056: begin
                        tc = f1055;
                        p1002 = p1002 - tc;
                        p983 = p983 + tc;
                end
                1057: begin
                        tc = f1056;
                        p140 = p140 - tc;
                        p1002 = p1002 + tc;
                end
                1058: begin
                        tc = f1057;
                        p1004 = p1004 - tc;
                        p1005 = p1005 + tc;
                end
                1059: begin
                        tc = f1058;
                        p1007 = p1007 - tc;
                        p1006 = p1006 + tc;
                end
                1060: begin
                        tc = f1059;
                        p146 = p146 - tc;
                        p1003 = p1003 + tc;
                        p1008 = p1008 + tc;
                end
                1061: begin
                        tc = f1060;
                        p1008 = p1008 - tc;
                        p146 = p146 + tc;
                end
                1062: begin
                        tc = f1061;
                        p1010 = p1010 - tc;
                        p1009 = p1009 + tc;
                end
                1063: begin
                        tc = f1062;
                        p1011 = p1011 - tc;
                        p1010 = p1010 + tc;
                end
                1064: begin
                        tc = f1063;
                        p149 = p149 - tc;
                        p1004 = p1004 + tc;
                        p1012 = p1012 + tc;
                end
                1065: begin
                        tc = f1064;
                        p1012 = p1012 - tc;
                        p149 = p149 + tc;
                end
                1066: begin
                        tc = f1065;
                        p1014 = p1014 - tc;
                        p1013 = p1013 + tc;
                end
                1067: begin
                        tc = f1066;
                        p1015 = p1015 - tc;
                        p1014 = p1014 + tc;
                end
                1068: begin
                        tc = f1067;
                        p1009 = p1009 - tc;
                        p1013 = p1013 - tc;
                        p140 = p140 + tc;
                end
                1069: begin
                        tc = f1068;
                        p1006 = p1006 - tc;
                        p1011 = p1011 + tc;
                        p1015 = p1015 + tc;
                end
                1070: begin
                        tc = f1069;
                        p1005 = p1005 - tc;
                        p150 = p150 + tc;
                end
                1071: begin
                        tc = f1070;
                        p150 = p150 - tc;
                end
                1072: begin
                        tc = f1071;
                        p1016 = p1016 - tc;
                        p1007 = p1007 + tc;
                end
                1073: begin
                        tc = f1072;
                        p141 = p141 - tc;
                        p1016 = p1016 + tc;
                end
                1074: begin
                        tc = f1073;
                        p1023 = p1023 - tc;
                        p1019 = p1019 + tc;
                end
                1075: begin
                        tc = f1074;
                        p1017 = p1017 - tc;
                end
                1076: begin
                        tc = f1075;
                        p1021 = p1021 - tc;
                        p1023 = p1023 + tc;
                end
                1077: begin
                        tc = f1076;
                        p1018 = p1018 - tc*2;
                        p1024 = p1024 + tc;
                end
                1078: begin
                        tc = f1077;
                        p1025 = p1025 - tc;
                        p1022 = p1022 + tc;
                end
                1079: begin
                        tc = f1078;
                        p1018 = p1018 - tc;
                        p1027 = p1027 - tc;
                        p1026 = p1026 + tc;
                end
                1080: begin
                        tc = f1079;
                        p1028 = p1028 - tc;
                        p1025 = p1025 + tc;
                end
                1081: begin
                        tc = f1080;
                        p1017 = p1017 - tc;
                        p1020 = p1020 + tc;
                        p1029 = p1029 + tc;
                end
                1082: begin
                        tc = f1081;
                        p1017 = p1017 - tc;
                        p1029 = p1029 + tc;
                end
                1083: begin
                        tc = f1082;
                        p1030 = p1030 - tc;
                        p1028 = p1028 + tc;
                end
                1084: begin
                        tc = f1083;
                        p1024 = p1024 - tc;
                        p1018 = p1018 + tc;
                end
                1085: begin
                        tc = f1084;
                        p1031 = p1031 - tc;
                        p1030 = p1030 + tc;
                end
                1086: begin
                        tc = f1085;
                        p1029 = p1029 - tc;
                        p1017 = p1017 + tc*2;
                end
                1087: begin
                        tc = f1086;
                        p1019 = p1019 - tc;
                        p1026 = p1026 - tc;
                        p1027 = p1027 + tc;
                        p1031 = p1031 + tc;
                end
                1088: begin
                        tc = f1087;
                        p1019 = p1019 - tc;
                        p1031 = p1031 + tc;
                end
                1089: begin
                        tc = f1088;
                        p151 = p151 - tc;
                        p1017 = p1017 + tc;
                        p1032 = p1032 + tc;
                end
                1090: begin
                        tc = f1089;
                        p1032 = p1032 - tc;
                        p151 = p151 + tc;
                end
                1091: begin
                        tc = f1090;
                        p1034 = p1034 - tc;
                        p1033 = p1033 + tc;
                end
                1092: begin
                        tc = f1091;
                        p1035 = p1035 - tc;
                        p1034 = p1034 + tc;
                end
                1093: begin
                        tc = f1092;
                        p152 = p152 - tc;
                        p1018 = p1018 + tc;
                        p1036 = p1036 + tc;
                end
                1094: begin
                        tc = f1093;
                        p1036 = p1036 - tc;
                        p152 = p152 + tc;
                end
                1095: begin
                        tc = f1094;
                        p1038 = p1038 - tc;
                        p1037 = p1037 + tc;
                end
                1096: begin
                        tc = f1095;
                        p1039 = p1039 - tc;
                        p1038 = p1038 + tc;
                end
                1097: begin
                        tc = f1096;
                        p1033 = p1033 - tc;
                        p1037 = p1037 - tc;
                        p141 = p141 + tc;
                end
                1098: begin
                        tc = f1097;
                        p1019 = p1019 - tc;
                        p1035 = p1035 + tc;
                        p1039 = p1039 + tc;
                end
                1099: begin
                        tc = f1098;
                        p1020 = p1020 - tc;
                        p153 = p153 + tc;
                end
                1100: begin
                        tc = f1099;
                        p153 = p153 - tc;
                end
                1101: begin
                        tc = f1100;
                        p1040 = p1040 - tc;
                        p1021 = p1021 + tc;
                end
                1102: begin
                        tc = f1101;
                        p142 = p142 - tc;
                        p1040 = p1040 + tc;
                end
                1103: begin
                        tc = f1102;
                        p1042 = p1042 - tc;
                        p1043 = p1043 + tc;
                end
                1104: begin
                        tc = f1103;
                        p1045 = p1045 - tc;
                        p1044 = p1044 + tc;
                end
                1105: begin
                        tc = f1104;
                        p150 = p150 - tc;
                        p1041 = p1041 + tc;
                        p1046 = p1046 + tc;
                end
                1106: begin
                        tc = f1105;
                        p1046 = p1046 - tc;
                        p150 = p150 + tc;
                end
                1107: begin
                        tc = f1106;
                        p1048 = p1048 - tc;
                        p1047 = p1047 + tc;
                end
                1108: begin
                        tc = f1107;
                        p1049 = p1049 - tc;
                        p1048 = p1048 + tc;
                end
                1109: begin
                        tc = f1108;
                        p153 = p153 - tc;
                        p1042 = p1042 + tc;
                        p1050 = p1050 + tc;
                end
                1110: begin
                        tc = f1109;
                        p1050 = p1050 - tc;
                        p153 = p153 + tc;
                end
                1111: begin
                        tc = f1110;
                        p1052 = p1052 - tc;
                        p1051 = p1051 + tc;
                end
                1112: begin
                        tc = f1111;
                        p1053 = p1053 - tc;
                        p1052 = p1052 + tc;
                end
                1113: begin
                        tc = f1112;
                        p1047 = p1047 - tc;
                        p1051 = p1051 - tc;
                        p142 = p142 + tc;
                end
                1114: begin
                        tc = f1113;
                        p1044 = p1044 - tc;
                        p1049 = p1049 + tc;
                        p1053 = p1053 + tc;
                end
                1115: begin
                        tc = f1114;
                        p1043 = p1043 - tc;
                        p154 = p154 + tc;
                end
                1116: begin
                        tc = f1115;
                        p154 = p154 - tc;
                end
                1117: begin
                        tc = f1116;
                        p1054 = p1054 - tc;
                        p1045 = p1045 + tc;
                end
                1118: begin
                        tc = f1117;
                        p143 = p143 - tc;
                        p1054 = p1054 + tc;
                end
                default:;
        endcase
        led = ~p18[5:0];
end
end
endmodule