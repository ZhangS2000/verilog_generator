module sn(
        input clk,
        output reg [5:0] led
);
`define INH(place) ((place) == 0 ? 2097151 : 0)
reg [20:0] p0=0,p1=1,p2=1,p3=1,p4=1,p5=1,p6=1,p7=1,p8=1,p9=1,p10=1,p11=1,p12=1,p13=1,p14=1,p15=8,p16=20,p17=0,p18=20,p19=0,p20=20,p21=0,p22=20,p23=0,p24=5,p25=20,p26=0,p27=20,p28=0,p29=20,p30=0,p31=0,p32=1,p33=20,p34=0,p35=20,p36=0,p37=0,p38=10,p39=20,p40=0,p41=0,p42=5,p43=0,p44=0,p45=0,p46=1,p47=0,p48=1,p49=1,p50=1,p51=0,p52=1,p53=0,p54=1,p55=1,p56=0,p57=1,p58=1,p59=0,p60=1,p61=1,p62=1,p63=0,p64=1,p65=1,p66=1,p67=1,p68=0,p69=0,p70=1,p71=0,p72=1,p73=1,p74=1,p75=0,p76=1,p77=0,p78=1,p79=1,p80=0,p81=1,p82=1,p83=0,p84=1,p85=1,p86=1,p87=0,p88=1,p89=1,p90=1,p91=1,p92=0,p93=0,p94=1,p95=0,p96=1,p97=1,p98=1,p99=0,p100=1,p101=0,p102=1,p103=1,p104=0,p105=1,p106=1,p107=0,p108=1,p109=1,p110=1,p111=0,p112=1,p113=1,p114=1,p115=1,p116=0,p117=0,p118=1,p119=0,p120=1,p121=1,p122=1,p123=0,p124=1,p125=0,p126=1,p127=1,p128=0,p129=1,p130=1,p131=0,p132=1,p133=1,p134=1,p135=0,p136=1,p137=1,p138=1,p139=1,p140=0,p141=0,p142=1,p143=0,p144=1,p145=1,p146=1,p147=0,p148=1,p149=0,p150=1,p151=1,p152=0,p153=1,p154=1,p155=0,p156=1,p157=1,p158=1,p159=0,p160=1,p161=1,p162=1,p163=1,p164=0,p165=0,p166=1,p167=0,p168=1,p169=1,p170=1,p171=0,p172=1,p173=0,p174=1,p175=1,p176=0,p177=1,p178=1,p179=0,p180=1,p181=1,p182=1,p183=0,p184=1,p185=1,p186=1,p187=1,p188=0,p189=0,p190=1,p191=0,p192=1,p193=1,p194=1,p195=0,p196=1,p197=0,p198=1,p199=1,p200=0,p201=1,p202=1,p203=0,p204=1,p205=1,p206=1,p207=0,p208=1,p209=1,p210=1,p211=1,p212=0,p213=0,p214=0,p215=1,p216=1,p217=0,p218=1,p219=1,p220=1,p221=0,p222=1,p223=1,p224=1,p225=1,p226=0,p227=0,p228=1,p229=0,p230=1,p231=1,p232=1,p233=0,p234=1,p235=0,p236=1,p237=1,p238=0,p239=1,p240=1,p241=0,p242=1,p243=1,p244=1,p245=0,p246=1,p247=1,p248=1,p249=1,p250=0,p251=0,p252=1,p253=0,p254=1,p255=1,p256=1,p257=0,p258=1,p259=0,p260=1,p261=1,p262=0,p263=1,p264=1,p265=0,p266=1,p267=1,p268=1,p269=0,p270=1,p271=1,p272=1,p273=1,p274=0,p275=0,p276=0,p277=1,p278=1,p279=0,p280=1,p281=1,p282=1,p283=0,p284=1,p285=1,p286=1,p287=1,p288=0,p289=0,p290=1,p291=0,p292=1,p293=1,p294=1,p295=0,p296=1,p297=0,p298=1,p299=1,p300=0,p301=1,p302=1,p303=0,p304=1,p305=1,p306=1,p307=0,p308=1,p309=1,p310=1,p311=1,p312=0,p313=0,p314=0,p315=1,p316=1,p317=0,p318=1,p319=1,p320=1,p321=0,p322=1,p323=1,p324=1,p325=1,p326=0,p327=0,p328=0,p329=1,p330=1,p331=0,p332=1,p333=1,p334=1,p335=0,p336=1,p337=1,p338=1,p339=1;
reg [20:0] f0,f1,f2,f3,f4,f5,f6,f7,f8,f9,f10,f11,f12,f13,f14,f15,f16,f17,f18,f19,f20,f21,f22,f23,f24,f25,f26,f27,f28,f29,f30,f31,f32,f33,f34,f35,f36,f37,f38,f39,f40,f41,f42,f43,f44,f45,f46,f47,f48,f49,f50,f51,f52,f53,f54,f55,f56,f57,f58,f59,f60,f61,f62,f63,f64,f65,f66,f67,f68,f69,f70,f71,f72,f73,f74,f75,f76,f77,f78,f79,f80,f81,f82,f83,f84,f85,f86,f87,f88,f89,f90,f91,f92,f93,f94,f95,f96,f97,f98,f99,f100,f101,f102,f103,f104,f105,f106,f107,f108,f109,f110,f111,f112,f113,f114,f115,f116,f117,f118,f119,f120,f121,f122,f123,f124,f125,f126,f127,f128,f129,f130,f131,f132,f133,f134,f135,f136,f137,f138,f139,f140,f141,f142,f143,f144,f145,f146,f147,f148,f149,f150,f151,f152,f153,f154,f155,f156,f157,f158,f159,f160,f161,f162,f163,f164,f165,f166,f167,f168,f169,f170,f171,f172,f173,f174,f175,f176,f177,f178,f179,f180,f181,f182,f183,f184,f185,f186,f187,f188,f189,f190,f191,f192,f193,f194,f195,f196,f197,f198,f199,f200,f201,f202,f203,f204,f205,f206,f207,f208,f209,f210,f211,f212,f213,f214,f215,f216,f217,f218,f219,f220,f221,f222,f223,f224,f225,f226,f227,f228,f229,f230,f231,f232,f233,f234,f235,f236,f237,f238,f239,f240,f241,f242,f243,f244,f245,f246,f247,f248,f249,f250,f251,f252,f253,f254,f255,f256,f257,f258,f259,f260,f261,f262,f263,f264,f265,f266,f267,f268,f269,f270,f271,f272,f273,f274,f275,f276,f277,f278,f279,f280,f281,f282,f283,f284,f285,f286,f287,f288,f289,f290,f291,f292,f293,f294,f295,f296,f297,f298,f299,f300,f301,f302,f303,f304,f305,f306,f307,f308,f309,f310,f311,f312,f313,f314,f315,f316,f317,f318,f319,f320,f321,f322,f323,f324,f325,f326,f327,f328,f329,f330,f331,f332,f333,f334,f335,f336,f337,f338,f339,f340,f341,f342,f343,f344,f345,f346,f347,f348,f349,f350,f351,f352,f353,f354,f355,f356,f357,f358,f359,f360,f361,f362,f363,f364,f365,f366,f367;
reg [20:0] tf;
reg [20:0] tc;
reg [47:0] counter1=1;
reg [1:0] clk_div; // 2位寄存器用于实现时钟分频

always @(posedge clk) begin
    if(clk_div < 2'b10)
        clk_div <= clk_div + 1; // 计数器自增
    else
        clk_div <= 2'b00; // 重置计数器
end

// 使用clk_div来控制某些逻辑的触发条件
always @(posedge clk) begin
    if (clk_div == 2'b10) begin
        f0 = 2097151;
        f0 = (f0 >= `INH(p46)) ? `INH(p46) : f0;
        f0 = (f0 > p49) ? p49 : f0;
        f1 = 2097151;
        f1 = (f1 >= `INH(p70)) ? `INH(p70) : f1;
        f1 = (f1 > p73) ? p73 : f1;
        f2 = 2097151;
        f2 = (f2 >= `INH(p94)) ? `INH(p94) : f2;
        f2 = (f2 > p97) ? p97 : f2;
        f3 = 2097151;
        f3 = (f3 >= `INH(p118)) ? `INH(p118) : f3;
        f3 = (f3 > p121) ? p121 : f3;
        f4 = 2097151;
        f4 = (f4 >= `INH(p142)) ? `INH(p142) : f4;
        f4 = (f4 > p145) ? p145 : f4;
        f5 = 2097151;
        f5 = (f5 >= `INH(p166)) ? `INH(p166) : f5;
        f5 = (f5 > p169) ? p169 : f5;
        f6 = 2097151;
        f6 = (f6 >= `INH(p190)) ? `INH(p190) : f6;
        f6 = (f6 > p193) ? p193 : f6;
        f7 = 2097151;
        f7 = (f7 > p212) ? p212 : f7;
        f7 = (f7 >= `INH(p215)) ? `INH(p215) : f7;
        f8 = 2097151;
        f8 = (f8 >= `INH(p228)) ? `INH(p228) : f8;
        f8 = (f8 > p231) ? p231 : f8;
        f9 = 2097151;
        f9 = (f9 >= `INH(p252)) ? `INH(p252) : f9;
        f9 = (f9 > p255) ? p255 : f9;
        f10 = 2097151;
        f10 = (f10 > p274) ? p274 : f10;
        f10 = (f10 >= `INH(p277)) ? `INH(p277) : f10;
        f11 = 2097151;
        f11 = (f11 >= `INH(p290)) ? `INH(p290) : f11;
        f11 = (f11 > p293) ? p293 : f11;
        f12 = 2097151;
        f12 = (f12 > p312) ? p312 : f12;
        f12 = (f12 >= `INH(p315)) ? `INH(p315) : f12;
        f13 = 2097151;
        f13 = (f13 > p326) ? p326 : f13;
        f13 = (f13 >= `INH(p329)) ? `INH(p329) : f13;
        f14 = 2097151;
        f14 = (f14 >= `INH(p45)) ? `INH(p45) : f14;
        f14 = (f14 >= `INH(p46)) ? `INH(p46) : f14;
        f14 = (f14 > p50) ? p50 : f14;
        f15 = 2097151;
        f15 = (f15 > p44) ? p44 : f15;
        f15 = (f15 >= `INH(p50)) ? `INH(p50) : f15;
        f16 = 2097151;
        f16 = (f16 > p48) ? p48 : f16;
        f16 = (f16 >= `INH(p50)) ? `INH(p50) : f16;
        f17 = 2097151;
        f17 = (f17 >= p45/2) ? p45/2 : f17;
        f17 = (f17 >= `INH(p49)) ? `INH(p49) : f17;
        f18 = 2097151;
        f18 = (f18 >= `INH(p49)) ? `INH(p49) : f18;
        f18 = (f18 > p52) ? p52 : f18;
        f19 = 2097151;
        f19 = (f19 > p45) ? p45 : f19;
        f19 = (f19 >= `INH(p52)) ? `INH(p52) : f19;
        f19 = (f19 > p54) ? p54 : f19;
        f20 = 2097151;
        f20 = (f20 >= `INH(p52)) ? `INH(p52) : f20;
        f20 = (f20 > p55) ? p55 : f20;
        f21 = 2097151;
        f21 = (f21 > p44) ? p44 : f21;
        f21 = (f21 >= `INH(p54)) ? `INH(p54) : f21;
        f21 = (f21 >= `INH(p55)) ? `INH(p55) : f21;
        f22 = 2097151;
        f22 = (f22 > p44) ? p44 : f22;
        f22 = (f22 >= `INH(p53)) ? `INH(p53) : f22;
        f22 = (f22 >= `INH(p55)) ? `INH(p55) : f22;
        f23 = 2097151;
        f23 = (f23 >= `INH(p55)) ? `INH(p55) : f23;
        f23 = (f23 > p57) ? p57 : f23;
        f24 = 2097151;
        f24 = (f24 > p51) ? p51 : f24;
        f24 = (f24 >= `INH(p57)) ? `INH(p57) : f24;
        f25 = 2097151;
        f25 = (f25 >= `INH(p57)) ? `INH(p57) : f25;
        f25 = (f25 > p58) ? p58 : f25;
        f26 = 2097151;
        f26 = (f26 > p56) ? p56 : f26;
        f26 = (f26 >= `INH(p58)) ? `INH(p58) : f26;
        f27 = 2097151;
        f27 = (f27 > p46) ? p46 : f27;
        f27 = (f27 > p53) ? p53 : f27;
        f27 = (f27 >= `INH(p54)) ? `INH(p54) : f27;
        f27 = (f27 >= `INH(p58)) ? `INH(p58) : f27;
        f28 = 2097151;
        f28 = (f28 > p46) ? p46 : f28;
        f28 = (f28 >= `INH(p53)) ? `INH(p53) : f28;
        f28 = (f28 >= `INH(p58)) ? `INH(p58) : f28;
        f29 = 2097151;
        f29 = (f29 > p15) ? p15 : f29;
        f29 = (f29 >= `INH(p60)) ? `INH(p60) : f29;
        f30 = 2097151;
        f30 = (f30 > p59) ? p59 : f30;
        f30 = (f30 >= `INH(p61)) ? `INH(p61) : f30;
        f31 = 2097151;
        f31 = (f31 >= `INH(p15)) ? `INH(p15) : f31;
        f31 = (f31 >= `INH(p60)) ? `INH(p60) : f31;
        f31 = (f31 > p61) ? p61 : f31;
        f32 = 2097151;
        f32 = (f32 >= `INH(p59)) ? `INH(p59) : f32;
        f32 = (f32 >= `INH(p61)) ? `INH(p61) : f32;
        f32 = (f32 > p62) ? p62 : f32;
        f33 = 2097151;
        f33 = (f33 > p16) ? p16 : f33;
        f33 = (f33 >= `INH(p64)) ? `INH(p64) : f33;
        f34 = 2097151;
        f34 = (f34 > p63) ? p63 : f34;
        f34 = (f34 >= `INH(p65)) ? `INH(p65) : f34;
        f35 = 2097151;
        f35 = (f35 >= `INH(p16)) ? `INH(p16) : f35;
        f35 = (f35 >= `INH(p64)) ? `INH(p64) : f35;
        f35 = (f35 > p65) ? p65 : f35;
        f36 = 2097151;
        f36 = (f36 >= `INH(p63)) ? `INH(p63) : f36;
        f36 = (f36 >= `INH(p65)) ? `INH(p65) : f36;
        f36 = (f36 > p66) ? p66 : f36;
        f37 = 2097151;
        f37 = (f37 >= `INH(p0)) ? `INH(p0) : f37;
        f37 = (f37 > p60) ? p60 : f37;
        f37 = (f37 > p64) ? p64 : f37;
        f38 = 2097151;
        f38 = (f38 > p46) ? p46 : f38;
        f38 = (f38 >= `INH(p62)) ? `INH(p62) : f38;
        f38 = (f38 >= `INH(p66)) ? `INH(p66) : f38;
        f39 = 2097151;
        f39 = (f39 > p47) ? p47 : f39;
        f39 = (f39 >= `INH(p67)) ? `INH(p67) : f39;
        f40 = 2097151;
        f40 = (f40 > p17) ? p17 : f40;
        f40 = (f40 >= `INH(p48)) ? `INH(p48) : f40;
        f41 = 2097151;
        f41 = (f41 >= `INH(p17)) ? `INH(p17) : f41;
        f41 = (f41 >= `INH(p48)) ? `INH(p48) : f41;
        f41 = (f41 > p67) ? p67 : f41;
        f42 = 2097151;
        f42 = (f42 > p1) ? p1 : f42;
        f42 = (f42 >= `INH(p47)) ? `INH(p47) : f42;
        f42 = (f42 >= `INH(p67)) ? `INH(p67) : f42;
        f43 = 2097151;
        f43 = (f43 >= `INH(p69)) ? `INH(p69) : f43;
        f43 = (f43 >= `INH(p70)) ? `INH(p70) : f43;
        f43 = (f43 > p74) ? p74 : f43;
        f44 = 2097151;
        f44 = (f44 > p68) ? p68 : f44;
        f44 = (f44 >= `INH(p74)) ? `INH(p74) : f44;
        f45 = 2097151;
        f45 = (f45 > p72) ? p72 : f45;
        f45 = (f45 >= `INH(p74)) ? `INH(p74) : f45;
        f46 = 2097151;
        f46 = (f46 >= p69/2) ? p69/2 : f46;
        f46 = (f46 >= `INH(p73)) ? `INH(p73) : f46;
        f47 = 2097151;
        f47 = (f47 >= `INH(p73)) ? `INH(p73) : f47;
        f47 = (f47 > p76) ? p76 : f47;
        f48 = 2097151;
        f48 = (f48 > p69) ? p69 : f48;
        f48 = (f48 >= `INH(p76)) ? `INH(p76) : f48;
        f48 = (f48 > p78) ? p78 : f48;
        f49 = 2097151;
        f49 = (f49 >= `INH(p76)) ? `INH(p76) : f49;
        f49 = (f49 > p79) ? p79 : f49;
        f50 = 2097151;
        f50 = (f50 > p68) ? p68 : f50;
        f50 = (f50 >= `INH(p78)) ? `INH(p78) : f50;
        f50 = (f50 >= `INH(p79)) ? `INH(p79) : f50;
        f51 = 2097151;
        f51 = (f51 > p68) ? p68 : f51;
        f51 = (f51 >= `INH(p77)) ? `INH(p77) : f51;
        f51 = (f51 >= `INH(p79)) ? `INH(p79) : f51;
        f52 = 2097151;
        f52 = (f52 >= `INH(p79)) ? `INH(p79) : f52;
        f52 = (f52 > p81) ? p81 : f52;
        f53 = 2097151;
        f53 = (f53 > p75) ? p75 : f53;
        f53 = (f53 >= `INH(p81)) ? `INH(p81) : f53;
        f54 = 2097151;
        f54 = (f54 >= `INH(p81)) ? `INH(p81) : f54;
        f54 = (f54 > p82) ? p82 : f54;
        f55 = 2097151;
        f55 = (f55 > p80) ? p80 : f55;
        f55 = (f55 >= `INH(p82)) ? `INH(p82) : f55;
        f56 = 2097151;
        f56 = (f56 > p70) ? p70 : f56;
        f56 = (f56 > p77) ? p77 : f56;
        f56 = (f56 >= `INH(p78)) ? `INH(p78) : f56;
        f56 = (f56 >= `INH(p82)) ? `INH(p82) : f56;
        f57 = 2097151;
        f57 = (f57 > p70) ? p70 : f57;
        f57 = (f57 >= `INH(p77)) ? `INH(p77) : f57;
        f57 = (f57 >= `INH(p82)) ? `INH(p82) : f57;
        f58 = 2097151;
        f58 = (f58 > p17) ? p17 : f58;
        f58 = (f58 >= `INH(p84)) ? `INH(p84) : f58;
        f59 = 2097151;
        f59 = (f59 > p83) ? p83 : f59;
        f59 = (f59 >= `INH(p85)) ? `INH(p85) : f59;
        f60 = 2097151;
        f60 = (f60 >= `INH(p17)) ? `INH(p17) : f60;
        f60 = (f60 >= `INH(p84)) ? `INH(p84) : f60;
        f60 = (f60 > p85) ? p85 : f60;
        f61 = 2097151;
        f61 = (f61 >= `INH(p83)) ? `INH(p83) : f61;
        f61 = (f61 >= `INH(p85)) ? `INH(p85) : f61;
        f61 = (f61 > p86) ? p86 : f61;
        f62 = 2097151;
        f62 = (f62 > p18) ? p18 : f62;
        f62 = (f62 >= `INH(p88)) ? `INH(p88) : f62;
        f63 = 2097151;
        f63 = (f63 > p87) ? p87 : f63;
        f63 = (f63 >= `INH(p89)) ? `INH(p89) : f63;
        f64 = 2097151;
        f64 = (f64 >= `INH(p18)) ? `INH(p18) : f64;
        f64 = (f64 >= `INH(p88)) ? `INH(p88) : f64;
        f64 = (f64 > p89) ? p89 : f64;
        f65 = 2097151;
        f65 = (f65 >= `INH(p87)) ? `INH(p87) : f65;
        f65 = (f65 >= `INH(p89)) ? `INH(p89) : f65;
        f65 = (f65 > p90) ? p90 : f65;
        f66 = 2097151;
        f66 = (f66 >= `INH(p1)) ? `INH(p1) : f66;
        f66 = (f66 > p84) ? p84 : f66;
        f66 = (f66 > p88) ? p88 : f66;
        f67 = 2097151;
        f67 = (f67 > p70) ? p70 : f67;
        f67 = (f67 >= `INH(p86)) ? `INH(p86) : f67;
        f67 = (f67 >= `INH(p90)) ? `INH(p90) : f67;
        f68 = 2097151;
        f68 = (f68 > p71) ? p71 : f68;
        f68 = (f68 >= `INH(p91)) ? `INH(p91) : f68;
        f69 = 2097151;
        f69 = (f69 > p19) ? p19 : f69;
        f69 = (f69 >= `INH(p72)) ? `INH(p72) : f69;
        f70 = 2097151;
        f70 = (f70 >= `INH(p19)) ? `INH(p19) : f70;
        f70 = (f70 >= `INH(p72)) ? `INH(p72) : f70;
        f70 = (f70 > p91) ? p91 : f70;
        f71 = 2097151;
        f71 = (f71 > p2) ? p2 : f71;
        f71 = (f71 >= `INH(p71)) ? `INH(p71) : f71;
        f71 = (f71 >= `INH(p91)) ? `INH(p91) : f71;
        f72 = 2097151;
        f72 = (f72 >= `INH(p93)) ? `INH(p93) : f72;
        f72 = (f72 >= `INH(p94)) ? `INH(p94) : f72;
        f72 = (f72 > p98) ? p98 : f72;
        f73 = 2097151;
        f73 = (f73 > p92) ? p92 : f73;
        f73 = (f73 >= `INH(p98)) ? `INH(p98) : f73;
        f74 = 2097151;
        f74 = (f74 > p96) ? p96 : f74;
        f74 = (f74 >= `INH(p98)) ? `INH(p98) : f74;
        f75 = 2097151;
        f75 = (f75 >= p93/2) ? p93/2 : f75;
        f75 = (f75 >= `INH(p97)) ? `INH(p97) : f75;
        f76 = 2097151;
        f76 = (f76 >= `INH(p97)) ? `INH(p97) : f76;
        f76 = (f76 > p100) ? p100 : f76;
        f77 = 2097151;
        f77 = (f77 > p93) ? p93 : f77;
        f77 = (f77 >= `INH(p100)) ? `INH(p100) : f77;
        f77 = (f77 > p102) ? p102 : f77;
        f78 = 2097151;
        f78 = (f78 >= `INH(p100)) ? `INH(p100) : f78;
        f78 = (f78 > p103) ? p103 : f78;
        f79 = 2097151;
        f79 = (f79 > p92) ? p92 : f79;
        f79 = (f79 >= `INH(p102)) ? `INH(p102) : f79;
        f79 = (f79 >= `INH(p103)) ? `INH(p103) : f79;
        f80 = 2097151;
        f80 = (f80 > p92) ? p92 : f80;
        f80 = (f80 >= `INH(p101)) ? `INH(p101) : f80;
        f80 = (f80 >= `INH(p103)) ? `INH(p103) : f80;
        f81 = 2097151;
        f81 = (f81 >= `INH(p103)) ? `INH(p103) : f81;
        f81 = (f81 > p105) ? p105 : f81;
        f82 = 2097151;
        f82 = (f82 > p99) ? p99 : f82;
        f82 = (f82 >= `INH(p105)) ? `INH(p105) : f82;
        f83 = 2097151;
        f83 = (f83 >= `INH(p105)) ? `INH(p105) : f83;
        f83 = (f83 > p106) ? p106 : f83;
        f84 = 2097151;
        f84 = (f84 > p104) ? p104 : f84;
        f84 = (f84 >= `INH(p106)) ? `INH(p106) : f84;
        f85 = 2097151;
        f85 = (f85 > p94) ? p94 : f85;
        f85 = (f85 > p101) ? p101 : f85;
        f85 = (f85 >= `INH(p102)) ? `INH(p102) : f85;
        f85 = (f85 >= `INH(p106)) ? `INH(p106) : f85;
        f86 = 2097151;
        f86 = (f86 > p94) ? p94 : f86;
        f86 = (f86 >= `INH(p101)) ? `INH(p101) : f86;
        f86 = (f86 >= `INH(p106)) ? `INH(p106) : f86;
        f87 = 2097151;
        f87 = (f87 > p19) ? p19 : f87;
        f87 = (f87 >= `INH(p108)) ? `INH(p108) : f87;
        f88 = 2097151;
        f88 = (f88 > p107) ? p107 : f88;
        f88 = (f88 >= `INH(p109)) ? `INH(p109) : f88;
        f89 = 2097151;
        f89 = (f89 >= `INH(p19)) ? `INH(p19) : f89;
        f89 = (f89 >= `INH(p108)) ? `INH(p108) : f89;
        f89 = (f89 > p109) ? p109 : f89;
        f90 = 2097151;
        f90 = (f90 >= `INH(p107)) ? `INH(p107) : f90;
        f90 = (f90 >= `INH(p109)) ? `INH(p109) : f90;
        f90 = (f90 > p110) ? p110 : f90;
        f91 = 2097151;
        f91 = (f91 > p20) ? p20 : f91;
        f91 = (f91 >= `INH(p112)) ? `INH(p112) : f91;
        f92 = 2097151;
        f92 = (f92 > p111) ? p111 : f92;
        f92 = (f92 >= `INH(p113)) ? `INH(p113) : f92;
        f93 = 2097151;
        f93 = (f93 >= `INH(p20)) ? `INH(p20) : f93;
        f93 = (f93 >= `INH(p112)) ? `INH(p112) : f93;
        f93 = (f93 > p113) ? p113 : f93;
        f94 = 2097151;
        f94 = (f94 >= `INH(p111)) ? `INH(p111) : f94;
        f94 = (f94 >= `INH(p113)) ? `INH(p113) : f94;
        f94 = (f94 > p114) ? p114 : f94;
        f95 = 2097151;
        f95 = (f95 >= `INH(p2)) ? `INH(p2) : f95;
        f95 = (f95 > p108) ? p108 : f95;
        f95 = (f95 > p112) ? p112 : f95;
        f96 = 2097151;
        f96 = (f96 > p94) ? p94 : f96;
        f96 = (f96 >= `INH(p110)) ? `INH(p110) : f96;
        f96 = (f96 >= `INH(p114)) ? `INH(p114) : f96;
        f97 = 2097151;
        f97 = (f97 > p95) ? p95 : f97;
        f97 = (f97 >= `INH(p115)) ? `INH(p115) : f97;
        f98 = 2097151;
        f98 = (f98 > p21) ? p21 : f98;
        f98 = (f98 >= `INH(p96)) ? `INH(p96) : f98;
        f99 = 2097151;
        f99 = (f99 >= `INH(p21)) ? `INH(p21) : f99;
        f99 = (f99 >= `INH(p96)) ? `INH(p96) : f99;
        f99 = (f99 > p115) ? p115 : f99;
        f100 = 2097151;
        f100 = (f100 > p3) ? p3 : f100;
        f100 = (f100 >= `INH(p95)) ? `INH(p95) : f100;
        f100 = (f100 >= `INH(p115)) ? `INH(p115) : f100;
        f101 = 2097151;
        f101 = (f101 >= `INH(p117)) ? `INH(p117) : f101;
        f101 = (f101 >= `INH(p118)) ? `INH(p118) : f101;
        f101 = (f101 > p122) ? p122 : f101;
        f102 = 2097151;
        f102 = (f102 > p116) ? p116 : f102;
        f102 = (f102 >= `INH(p122)) ? `INH(p122) : f102;
        f103 = 2097151;
        f103 = (f103 > p120) ? p120 : f103;
        f103 = (f103 >= `INH(p122)) ? `INH(p122) : f103;
        f104 = 2097151;
        f104 = (f104 >= p117/2) ? p117/2 : f104;
        f104 = (f104 >= `INH(p121)) ? `INH(p121) : f104;
        f105 = 2097151;
        f105 = (f105 >= `INH(p121)) ? `INH(p121) : f105;
        f105 = (f105 > p124) ? p124 : f105;
        f106 = 2097151;
        f106 = (f106 > p117) ? p117 : f106;
        f106 = (f106 >= `INH(p124)) ? `INH(p124) : f106;
        f106 = (f106 > p126) ? p126 : f106;
        f107 = 2097151;
        f107 = (f107 >= `INH(p124)) ? `INH(p124) : f107;
        f107 = (f107 > p127) ? p127 : f107;
        f108 = 2097151;
        f108 = (f108 > p116) ? p116 : f108;
        f108 = (f108 >= `INH(p126)) ? `INH(p126) : f108;
        f108 = (f108 >= `INH(p127)) ? `INH(p127) : f108;
        f109 = 2097151;
        f109 = (f109 > p116) ? p116 : f109;
        f109 = (f109 >= `INH(p125)) ? `INH(p125) : f109;
        f109 = (f109 >= `INH(p127)) ? `INH(p127) : f109;
        f110 = 2097151;
        f110 = (f110 >= `INH(p127)) ? `INH(p127) : f110;
        f110 = (f110 > p129) ? p129 : f110;
        f111 = 2097151;
        f111 = (f111 > p123) ? p123 : f111;
        f111 = (f111 >= `INH(p129)) ? `INH(p129) : f111;
        f112 = 2097151;
        f112 = (f112 >= `INH(p129)) ? `INH(p129) : f112;
        f112 = (f112 > p130) ? p130 : f112;
        f113 = 2097151;
        f113 = (f113 > p128) ? p128 : f113;
        f113 = (f113 >= `INH(p130)) ? `INH(p130) : f113;
        f114 = 2097151;
        f114 = (f114 > p118) ? p118 : f114;
        f114 = (f114 > p125) ? p125 : f114;
        f114 = (f114 >= `INH(p126)) ? `INH(p126) : f114;
        f114 = (f114 >= `INH(p130)) ? `INH(p130) : f114;
        f115 = 2097151;
        f115 = (f115 > p118) ? p118 : f115;
        f115 = (f115 >= `INH(p125)) ? `INH(p125) : f115;
        f115 = (f115 >= `INH(p130)) ? `INH(p130) : f115;
        f116 = 2097151;
        f116 = (f116 > p21) ? p21 : f116;
        f116 = (f116 >= `INH(p132)) ? `INH(p132) : f116;
        f117 = 2097151;
        f117 = (f117 > p131) ? p131 : f117;
        f117 = (f117 >= `INH(p133)) ? `INH(p133) : f117;
        f118 = 2097151;
        f118 = (f118 >= `INH(p21)) ? `INH(p21) : f118;
        f118 = (f118 >= `INH(p132)) ? `INH(p132) : f118;
        f118 = (f118 > p133) ? p133 : f118;
        f119 = 2097151;
        f119 = (f119 >= `INH(p131)) ? `INH(p131) : f119;
        f119 = (f119 >= `INH(p133)) ? `INH(p133) : f119;
        f119 = (f119 > p134) ? p134 : f119;
        f120 = 2097151;
        f120 = (f120 > p22) ? p22 : f120;
        f120 = (f120 >= `INH(p136)) ? `INH(p136) : f120;
        f121 = 2097151;
        f121 = (f121 > p135) ? p135 : f121;
        f121 = (f121 >= `INH(p137)) ? `INH(p137) : f121;
        f122 = 2097151;
        f122 = (f122 >= `INH(p22)) ? `INH(p22) : f122;
        f122 = (f122 >= `INH(p136)) ? `INH(p136) : f122;
        f122 = (f122 > p137) ? p137 : f122;
        f123 = 2097151;
        f123 = (f123 >= `INH(p135)) ? `INH(p135) : f123;
        f123 = (f123 >= `INH(p137)) ? `INH(p137) : f123;
        f123 = (f123 > p138) ? p138 : f123;
        f124 = 2097151;
        f124 = (f124 >= `INH(p3)) ? `INH(p3) : f124;
        f124 = (f124 > p132) ? p132 : f124;
        f124 = (f124 > p136) ? p136 : f124;
        f125 = 2097151;
        f125 = (f125 > p118) ? p118 : f125;
        f125 = (f125 >= `INH(p134)) ? `INH(p134) : f125;
        f125 = (f125 >= `INH(p138)) ? `INH(p138) : f125;
        f126 = 2097151;
        f126 = (f126 > p119) ? p119 : f126;
        f126 = (f126 >= `INH(p139)) ? `INH(p139) : f126;
        f127 = 2097151;
        f127 = (f127 > p23) ? p23 : f127;
        f127 = (f127 >= `INH(p120)) ? `INH(p120) : f127;
        f128 = 2097151;
        f128 = (f128 >= `INH(p23)) ? `INH(p23) : f128;
        f128 = (f128 >= `INH(p120)) ? `INH(p120) : f128;
        f128 = (f128 > p139) ? p139 : f128;
        f129 = 2097151;
        f129 = (f129 > p4) ? p4 : f129;
        f129 = (f129 >= `INH(p119)) ? `INH(p119) : f129;
        f129 = (f129 >= `INH(p139)) ? `INH(p139) : f129;
        f130 = 2097151;
        f130 = (f130 >= `INH(p141)) ? `INH(p141) : f130;
        f130 = (f130 >= `INH(p142)) ? `INH(p142) : f130;
        f130 = (f130 > p146) ? p146 : f130;
        f131 = 2097151;
        f131 = (f131 > p140) ? p140 : f131;
        f131 = (f131 >= `INH(p146)) ? `INH(p146) : f131;
        f132 = 2097151;
        f132 = (f132 > p144) ? p144 : f132;
        f132 = (f132 >= `INH(p146)) ? `INH(p146) : f132;
        f133 = 2097151;
        f133 = (f133 >= p141/2) ? p141/2 : f133;
        f133 = (f133 >= `INH(p145)) ? `INH(p145) : f133;
        f134 = 2097151;
        f134 = (f134 >= `INH(p145)) ? `INH(p145) : f134;
        f134 = (f134 > p148) ? p148 : f134;
        f135 = 2097151;
        f135 = (f135 > p141) ? p141 : f135;
        f135 = (f135 >= `INH(p148)) ? `INH(p148) : f135;
        f135 = (f135 > p150) ? p150 : f135;
        f136 = 2097151;
        f136 = (f136 >= `INH(p148)) ? `INH(p148) : f136;
        f136 = (f136 > p151) ? p151 : f136;
        f137 = 2097151;
        f137 = (f137 > p140) ? p140 : f137;
        f137 = (f137 >= `INH(p150)) ? `INH(p150) : f137;
        f137 = (f137 >= `INH(p151)) ? `INH(p151) : f137;
        f138 = 2097151;
        f138 = (f138 > p140) ? p140 : f138;
        f138 = (f138 >= `INH(p149)) ? `INH(p149) : f138;
        f138 = (f138 >= `INH(p151)) ? `INH(p151) : f138;
        f139 = 2097151;
        f139 = (f139 >= `INH(p151)) ? `INH(p151) : f139;
        f139 = (f139 > p153) ? p153 : f139;
        f140 = 2097151;
        f140 = (f140 > p147) ? p147 : f140;
        f140 = (f140 >= `INH(p153)) ? `INH(p153) : f140;
        f141 = 2097151;
        f141 = (f141 >= `INH(p153)) ? `INH(p153) : f141;
        f141 = (f141 > p154) ? p154 : f141;
        f142 = 2097151;
        f142 = (f142 > p152) ? p152 : f142;
        f142 = (f142 >= `INH(p154)) ? `INH(p154) : f142;
        f143 = 2097151;
        f143 = (f143 > p142) ? p142 : f143;
        f143 = (f143 > p149) ? p149 : f143;
        f143 = (f143 >= `INH(p150)) ? `INH(p150) : f143;
        f143 = (f143 >= `INH(p154)) ? `INH(p154) : f143;
        f144 = 2097151;
        f144 = (f144 > p142) ? p142 : f144;
        f144 = (f144 >= `INH(p149)) ? `INH(p149) : f144;
        f144 = (f144 >= `INH(p154)) ? `INH(p154) : f144;
        f145 = 2097151;
        f145 = (f145 > p24) ? p24 : f145;
        f145 = (f145 >= `INH(p156)) ? `INH(p156) : f145;
        f146 = 2097151;
        f146 = (f146 > p155) ? p155 : f146;
        f146 = (f146 >= `INH(p157)) ? `INH(p157) : f146;
        f147 = 2097151;
        f147 = (f147 >= `INH(p24)) ? `INH(p24) : f147;
        f147 = (f147 >= `INH(p156)) ? `INH(p156) : f147;
        f147 = (f147 > p157) ? p157 : f147;
        f148 = 2097151;
        f148 = (f148 >= `INH(p155)) ? `INH(p155) : f148;
        f148 = (f148 >= `INH(p157)) ? `INH(p157) : f148;
        f148 = (f148 > p158) ? p158 : f148;
        f149 = 2097151;
        f149 = (f149 > p25) ? p25 : f149;
        f149 = (f149 >= `INH(p160)) ? `INH(p160) : f149;
        f150 = 2097151;
        f150 = (f150 > p159) ? p159 : f150;
        f150 = (f150 >= `INH(p161)) ? `INH(p161) : f150;
        f151 = 2097151;
        f151 = (f151 >= `INH(p25)) ? `INH(p25) : f151;
        f151 = (f151 >= `INH(p160)) ? `INH(p160) : f151;
        f151 = (f151 > p161) ? p161 : f151;
        f152 = 2097151;
        f152 = (f152 >= `INH(p159)) ? `INH(p159) : f152;
        f152 = (f152 >= `INH(p161)) ? `INH(p161) : f152;
        f152 = (f152 > p162) ? p162 : f152;
        f153 = 2097151;
        f153 = (f153 >= `INH(p4)) ? `INH(p4) : f153;
        f153 = (f153 > p156) ? p156 : f153;
        f153 = (f153 > p160) ? p160 : f153;
        f154 = 2097151;
        f154 = (f154 > p142) ? p142 : f154;
        f154 = (f154 >= `INH(p158)) ? `INH(p158) : f154;
        f154 = (f154 >= `INH(p162)) ? `INH(p162) : f154;
        f155 = 2097151;
        f155 = (f155 > p143) ? p143 : f155;
        f155 = (f155 >= `INH(p163)) ? `INH(p163) : f155;
        f156 = 2097151;
        f156 = (f156 > p26) ? p26 : f156;
        f156 = (f156 >= `INH(p144)) ? `INH(p144) : f156;
        f157 = 2097151;
        f157 = (f157 >= `INH(p26)) ? `INH(p26) : f157;
        f157 = (f157 >= `INH(p144)) ? `INH(p144) : f157;
        f157 = (f157 > p163) ? p163 : f157;
        f158 = 2097151;
        f158 = (f158 > p5) ? p5 : f158;
        f158 = (f158 >= `INH(p143)) ? `INH(p143) : f158;
        f158 = (f158 >= `INH(p163)) ? `INH(p163) : f158;
        f159 = 2097151;
        f159 = (f159 >= `INH(p165)) ? `INH(p165) : f159;
        f159 = (f159 >= `INH(p166)) ? `INH(p166) : f159;
        f159 = (f159 > p170) ? p170 : f159;
        f160 = 2097151;
        f160 = (f160 > p164) ? p164 : f160;
        f160 = (f160 >= `INH(p170)) ? `INH(p170) : f160;
        f161 = 2097151;
        f161 = (f161 > p168) ? p168 : f161;
        f161 = (f161 >= `INH(p170)) ? `INH(p170) : f161;
        f162 = 2097151;
        f162 = (f162 >= p165/2) ? p165/2 : f162;
        f162 = (f162 >= `INH(p169)) ? `INH(p169) : f162;
        f163 = 2097151;
        f163 = (f163 >= `INH(p169)) ? `INH(p169) : f163;
        f163 = (f163 > p172) ? p172 : f163;
        f164 = 2097151;
        f164 = (f164 > p165) ? p165 : f164;
        f164 = (f164 >= `INH(p172)) ? `INH(p172) : f164;
        f164 = (f164 > p174) ? p174 : f164;
        f165 = 2097151;
        f165 = (f165 >= `INH(p172)) ? `INH(p172) : f165;
        f165 = (f165 > p175) ? p175 : f165;
        f166 = 2097151;
        f166 = (f166 > p164) ? p164 : f166;
        f166 = (f166 >= `INH(p174)) ? `INH(p174) : f166;
        f166 = (f166 >= `INH(p175)) ? `INH(p175) : f166;
        f167 = 2097151;
        f167 = (f167 > p164) ? p164 : f167;
        f167 = (f167 >= `INH(p173)) ? `INH(p173) : f167;
        f167 = (f167 >= `INH(p175)) ? `INH(p175) : f167;
        f168 = 2097151;
        f168 = (f168 >= `INH(p175)) ? `INH(p175) : f168;
        f168 = (f168 > p177) ? p177 : f168;
        f169 = 2097151;
        f169 = (f169 > p171) ? p171 : f169;
        f169 = (f169 >= `INH(p177)) ? `INH(p177) : f169;
        f170 = 2097151;
        f170 = (f170 >= `INH(p177)) ? `INH(p177) : f170;
        f170 = (f170 > p178) ? p178 : f170;
        f171 = 2097151;
        f171 = (f171 > p176) ? p176 : f171;
        f171 = (f171 >= `INH(p178)) ? `INH(p178) : f171;
        f172 = 2097151;
        f172 = (f172 > p166) ? p166 : f172;
        f172 = (f172 > p173) ? p173 : f172;
        f172 = (f172 >= `INH(p174)) ? `INH(p174) : f172;
        f172 = (f172 >= `INH(p178)) ? `INH(p178) : f172;
        f173 = 2097151;
        f173 = (f173 > p166) ? p166 : f173;
        f173 = (f173 >= `INH(p173)) ? `INH(p173) : f173;
        f173 = (f173 >= `INH(p178)) ? `INH(p178) : f173;
        f174 = 2097151;
        f174 = (f174 > p26) ? p26 : f174;
        f174 = (f174 >= `INH(p180)) ? `INH(p180) : f174;
        f175 = 2097151;
        f175 = (f175 > p179) ? p179 : f175;
        f175 = (f175 >= `INH(p181)) ? `INH(p181) : f175;
        f176 = 2097151;
        f176 = (f176 >= `INH(p26)) ? `INH(p26) : f176;
        f176 = (f176 >= `INH(p180)) ? `INH(p180) : f176;
        f176 = (f176 > p181) ? p181 : f176;
        f177 = 2097151;
        f177 = (f177 >= `INH(p179)) ? `INH(p179) : f177;
        f177 = (f177 >= `INH(p181)) ? `INH(p181) : f177;
        f177 = (f177 > p182) ? p182 : f177;
        f178 = 2097151;
        f178 = (f178 > p27) ? p27 : f178;
        f178 = (f178 >= `INH(p184)) ? `INH(p184) : f178;
        f179 = 2097151;
        f179 = (f179 > p183) ? p183 : f179;
        f179 = (f179 >= `INH(p185)) ? `INH(p185) : f179;
        f180 = 2097151;
        f180 = (f180 >= `INH(p27)) ? `INH(p27) : f180;
        f180 = (f180 >= `INH(p184)) ? `INH(p184) : f180;
        f180 = (f180 > p185) ? p185 : f180;
        f181 = 2097151;
        f181 = (f181 >= `INH(p183)) ? `INH(p183) : f181;
        f181 = (f181 >= `INH(p185)) ? `INH(p185) : f181;
        f181 = (f181 > p186) ? p186 : f181;
        f182 = 2097151;
        f182 = (f182 >= `INH(p5)) ? `INH(p5) : f182;
        f182 = (f182 > p180) ? p180 : f182;
        f182 = (f182 > p184) ? p184 : f182;
        f183 = 2097151;
        f183 = (f183 > p166) ? p166 : f183;
        f183 = (f183 >= `INH(p182)) ? `INH(p182) : f183;
        f183 = (f183 >= `INH(p186)) ? `INH(p186) : f183;
        f184 = 2097151;
        f184 = (f184 > p167) ? p167 : f184;
        f184 = (f184 >= `INH(p187)) ? `INH(p187) : f184;
        f185 = 2097151;
        f185 = (f185 > p28) ? p28 : f185;
        f185 = (f185 >= `INH(p168)) ? `INH(p168) : f185;
        f186 = 2097151;
        f186 = (f186 >= `INH(p28)) ? `INH(p28) : f186;
        f186 = (f186 >= `INH(p168)) ? `INH(p168) : f186;
        f186 = (f186 > p187) ? p187 : f186;
        f187 = 2097151;
        f187 = (f187 > p6) ? p6 : f187;
        f187 = (f187 >= `INH(p167)) ? `INH(p167) : f187;
        f187 = (f187 >= `INH(p187)) ? `INH(p187) : f187;
        f188 = 2097151;
        f188 = (f188 >= `INH(p189)) ? `INH(p189) : f188;
        f188 = (f188 >= `INH(p190)) ? `INH(p190) : f188;
        f188 = (f188 > p194) ? p194 : f188;
        f189 = 2097151;
        f189 = (f189 > p188) ? p188 : f189;
        f189 = (f189 >= `INH(p194)) ? `INH(p194) : f189;
        f190 = 2097151;
        f190 = (f190 > p192) ? p192 : f190;
        f190 = (f190 >= `INH(p194)) ? `INH(p194) : f190;
        f191 = 2097151;
        f191 = (f191 >= p189/2) ? p189/2 : f191;
        f191 = (f191 >= `INH(p193)) ? `INH(p193) : f191;
        f192 = 2097151;
        f192 = (f192 >= `INH(p193)) ? `INH(p193) : f192;
        f192 = (f192 > p196) ? p196 : f192;
        f193 = 2097151;
        f193 = (f193 > p189) ? p189 : f193;
        f193 = (f193 >= `INH(p196)) ? `INH(p196) : f193;
        f193 = (f193 > p198) ? p198 : f193;
        f194 = 2097151;
        f194 = (f194 >= `INH(p196)) ? `INH(p196) : f194;
        f194 = (f194 > p199) ? p199 : f194;
        f195 = 2097151;
        f195 = (f195 > p188) ? p188 : f195;
        f195 = (f195 >= `INH(p198)) ? `INH(p198) : f195;
        f195 = (f195 >= `INH(p199)) ? `INH(p199) : f195;
        f196 = 2097151;
        f196 = (f196 > p188) ? p188 : f196;
        f196 = (f196 >= `INH(p197)) ? `INH(p197) : f196;
        f196 = (f196 >= `INH(p199)) ? `INH(p199) : f196;
        f197 = 2097151;
        f197 = (f197 >= `INH(p199)) ? `INH(p199) : f197;
        f197 = (f197 > p201) ? p201 : f197;
        f198 = 2097151;
        f198 = (f198 > p195) ? p195 : f198;
        f198 = (f198 >= `INH(p201)) ? `INH(p201) : f198;
        f199 = 2097151;
        f199 = (f199 >= `INH(p201)) ? `INH(p201) : f199;
        f199 = (f199 > p202) ? p202 : f199;
        f200 = 2097151;
        f200 = (f200 > p200) ? p200 : f200;
        f200 = (f200 >= `INH(p202)) ? `INH(p202) : f200;
        f201 = 2097151;
        f201 = (f201 > p190) ? p190 : f201;
        f201 = (f201 > p197) ? p197 : f201;
        f201 = (f201 >= `INH(p198)) ? `INH(p198) : f201;
        f201 = (f201 >= `INH(p202)) ? `INH(p202) : f201;
        f202 = 2097151;
        f202 = (f202 > p190) ? p190 : f202;
        f202 = (f202 >= `INH(p197)) ? `INH(p197) : f202;
        f202 = (f202 >= `INH(p202)) ? `INH(p202) : f202;
        f203 = 2097151;
        f203 = (f203 > p28) ? p28 : f203;
        f203 = (f203 >= `INH(p204)) ? `INH(p204) : f203;
        f204 = 2097151;
        f204 = (f204 > p203) ? p203 : f204;
        f204 = (f204 >= `INH(p205)) ? `INH(p205) : f204;
        f205 = 2097151;
        f205 = (f205 >= `INH(p28)) ? `INH(p28) : f205;
        f205 = (f205 >= `INH(p204)) ? `INH(p204) : f205;
        f205 = (f205 > p205) ? p205 : f205;
        f206 = 2097151;
        f206 = (f206 >= `INH(p203)) ? `INH(p203) : f206;
        f206 = (f206 >= `INH(p205)) ? `INH(p205) : f206;
        f206 = (f206 > p206) ? p206 : f206;
        f207 = 2097151;
        f207 = (f207 > p29) ? p29 : f207;
        f207 = (f207 >= `INH(p208)) ? `INH(p208) : f207;
        f208 = 2097151;
        f208 = (f208 > p207) ? p207 : f208;
        f208 = (f208 >= `INH(p209)) ? `INH(p209) : f208;
        f209 = 2097151;
        f209 = (f209 >= `INH(p29)) ? `INH(p29) : f209;
        f209 = (f209 >= `INH(p208)) ? `INH(p208) : f209;
        f209 = (f209 > p209) ? p209 : f209;
        f210 = 2097151;
        f210 = (f210 >= `INH(p207)) ? `INH(p207) : f210;
        f210 = (f210 >= `INH(p209)) ? `INH(p209) : f210;
        f210 = (f210 > p210) ? p210 : f210;
        f211 = 2097151;
        f211 = (f211 >= `INH(p6)) ? `INH(p6) : f211;
        f211 = (f211 > p204) ? p204 : f211;
        f211 = (f211 > p208) ? p208 : f211;
        f212 = 2097151;
        f212 = (f212 > p190) ? p190 : f212;
        f212 = (f212 >= `INH(p206)) ? `INH(p206) : f212;
        f212 = (f212 >= `INH(p210)) ? `INH(p210) : f212;
        f213 = 2097151;
        f213 = (f213 > p191) ? p191 : f213;
        f213 = (f213 >= `INH(p211)) ? `INH(p211) : f213;
        f214 = 2097151;
        f214 = (f214 > p30) ? p30 : f214;
        f214 = (f214 >= `INH(p192)) ? `INH(p192) : f214;
        f215 = 2097151;
        f215 = (f215 >= `INH(p30)) ? `INH(p30) : f215;
        f215 = (f215 >= `INH(p192)) ? `INH(p192) : f215;
        f215 = (f215 > p211) ? p211 : f215;
        f216 = 2097151;
        f216 = (f216 > p7) ? p7 : f216;
        f216 = (f216 >= `INH(p191)) ? `INH(p191) : f216;
        f216 = (f216 >= `INH(p211)) ? `INH(p211) : f216;
        f217 = 2097151;
        f217 = (f217 > p213) ? p213 : f217;
        f217 = (f217 >= `INH(p215)) ? `INH(p215) : f217;
        f218 = 2097151;
        f218 = (f218 >= `INH(p212)) ? `INH(p212) : f218;
        f218 = (f218 >= `INH(p213)) ? `INH(p213) : f218;
        f218 = (f218 >= `INH(p215)) ? `INH(p215) : f218;
        f218 = (f218 > p216) ? p216 : f218;
        f219 = 2097151;
        f219 = (f219 > p23) ? p23 : f219;
        f219 = (f219 >= `INH(p218)) ? `INH(p218) : f219;
        f220 = 2097151;
        f220 = (f220 > p217) ? p217 : f220;
        f220 = (f220 >= `INH(p219)) ? `INH(p219) : f220;
        f221 = 2097151;
        f221 = (f221 >= `INH(p23)) ? `INH(p23) : f221;
        f221 = (f221 >= `INH(p218)) ? `INH(p218) : f221;
        f221 = (f221 > p219) ? p219 : f221;
        f222 = 2097151;
        f222 = (f222 >= `INH(p217)) ? `INH(p217) : f222;
        f222 = (f222 >= `INH(p219)) ? `INH(p219) : f222;
        f222 = (f222 > p220) ? p220 : f222;
        f223 = 2097151;
        f223 = (f223 > p30) ? p30 : f223;
        f223 = (f223 >= `INH(p222)) ? `INH(p222) : f223;
        f224 = 2097151;
        f224 = (f224 > p221) ? p221 : f224;
        f224 = (f224 >= `INH(p223)) ? `INH(p223) : f224;
        f225 = 2097151;
        f225 = (f225 >= `INH(p30)) ? `INH(p30) : f225;
        f225 = (f225 >= `INH(p222)) ? `INH(p222) : f225;
        f225 = (f225 > p223) ? p223 : f225;
        f226 = 2097151;
        f226 = (f226 >= `INH(p221)) ? `INH(p221) : f226;
        f226 = (f226 >= `INH(p223)) ? `INH(p223) : f226;
        f226 = (f226 > p224) ? p224 : f226;
        f227 = 2097151;
        f227 = (f227 >= `INH(p7)) ? `INH(p7) : f227;
        f227 = (f227 > p218) ? p218 : f227;
        f227 = (f227 > p222) ? p222 : f227;
        f228 = 2097151;
        f228 = (f228 > p215) ? p215 : f228;
        f228 = (f228 >= `INH(p220)) ? `INH(p220) : f228;
        f228 = (f228 >= `INH(p224)) ? `INH(p224) : f228;
        f229 = 2097151;
        f229 = (f229 > p214) ? p214 : f229;
        f229 = (f229 >= `INH(p225)) ? `INH(p225) : f229;
        f230 = 2097151;
        f230 = (f230 > p31) ? p31 : f230;
        f230 = (f230 >= `INH(p216)) ? `INH(p216) : f230;
        f231 = 2097151;
        f231 = (f231 >= `INH(p31)) ? `INH(p31) : f231;
        f231 = (f231 >= `INH(p216)) ? `INH(p216) : f231;
        f231 = (f231 > p225) ? p225 : f231;
        f232 = 2097151;
        f232 = (f232 > p8) ? p8 : f232;
        f232 = (f232 >= `INH(p214)) ? `INH(p214) : f232;
        f232 = (f232 >= `INH(p225)) ? `INH(p225) : f232;
        f233 = 2097151;
        f233 = (f233 >= `INH(p227)) ? `INH(p227) : f233;
        f233 = (f233 >= `INH(p228)) ? `INH(p228) : f233;
        f233 = (f233 > p232) ? p232 : f233;
        f234 = 2097151;
        f234 = (f234 > p226) ? p226 : f234;
        f234 = (f234 >= `INH(p232)) ? `INH(p232) : f234;
        f235 = 2097151;
        f235 = (f235 > p230) ? p230 : f235;
        f235 = (f235 >= `INH(p232)) ? `INH(p232) : f235;
        f236 = 2097151;
        f236 = (f236 >= p227/2) ? p227/2 : f236;
        f236 = (f236 >= `INH(p231)) ? `INH(p231) : f236;
        f237 = 2097151;
        f237 = (f237 >= `INH(p231)) ? `INH(p231) : f237;
        f237 = (f237 > p234) ? p234 : f237;
        f238 = 2097151;
        f238 = (f238 > p227) ? p227 : f238;
        f238 = (f238 >= `INH(p234)) ? `INH(p234) : f238;
        f238 = (f238 > p236) ? p236 : f238;
        f239 = 2097151;
        f239 = (f239 >= `INH(p234)) ? `INH(p234) : f239;
        f239 = (f239 > p237) ? p237 : f239;
        f240 = 2097151;
        f240 = (f240 > p226) ? p226 : f240;
        f240 = (f240 >= `INH(p236)) ? `INH(p236) : f240;
        f240 = (f240 >= `INH(p237)) ? `INH(p237) : f240;
        f241 = 2097151;
        f241 = (f241 > p226) ? p226 : f241;
        f241 = (f241 >= `INH(p235)) ? `INH(p235) : f241;
        f241 = (f241 >= `INH(p237)) ? `INH(p237) : f241;
        f242 = 2097151;
        f242 = (f242 >= `INH(p237)) ? `INH(p237) : f242;
        f242 = (f242 > p239) ? p239 : f242;
        f243 = 2097151;
        f243 = (f243 > p233) ? p233 : f243;
        f243 = (f243 >= `INH(p239)) ? `INH(p239) : f243;
        f244 = 2097151;
        f244 = (f244 >= `INH(p239)) ? `INH(p239) : f244;
        f244 = (f244 > p240) ? p240 : f244;
        f245 = 2097151;
        f245 = (f245 > p238) ? p238 : f245;
        f245 = (f245 >= `INH(p240)) ? `INH(p240) : f245;
        f246 = 2097151;
        f246 = (f246 > p228) ? p228 : f246;
        f246 = (f246 > p235) ? p235 : f246;
        f246 = (f246 >= `INH(p236)) ? `INH(p236) : f246;
        f246 = (f246 >= `INH(p240)) ? `INH(p240) : f246;
        f247 = 2097151;
        f247 = (f247 > p228) ? p228 : f247;
        f247 = (f247 >= `INH(p235)) ? `INH(p235) : f247;
        f247 = (f247 >= `INH(p240)) ? `INH(p240) : f247;
        f248 = 2097151;
        f248 = (f248 > p32) ? p32 : f248;
        f248 = (f248 >= `INH(p242)) ? `INH(p242) : f248;
        f249 = 2097151;
        f249 = (f249 > p241) ? p241 : f249;
        f249 = (f249 >= `INH(p243)) ? `INH(p243) : f249;
        f250 = 2097151;
        f250 = (f250 >= `INH(p32)) ? `INH(p32) : f250;
        f250 = (f250 >= `INH(p242)) ? `INH(p242) : f250;
        f250 = (f250 > p243) ? p243 : f250;
        f251 = 2097151;
        f251 = (f251 >= `INH(p241)) ? `INH(p241) : f251;
        f251 = (f251 >= `INH(p243)) ? `INH(p243) : f251;
        f251 = (f251 > p244) ? p244 : f251;
        f252 = 2097151;
        f252 = (f252 > p33) ? p33 : f252;
        f252 = (f252 >= `INH(p246)) ? `INH(p246) : f252;
        f253 = 2097151;
        f253 = (f253 > p245) ? p245 : f253;
        f253 = (f253 >= `INH(p247)) ? `INH(p247) : f253;
        f254 = 2097151;
        f254 = (f254 >= `INH(p33)) ? `INH(p33) : f254;
        f254 = (f254 >= `INH(p246)) ? `INH(p246) : f254;
        f254 = (f254 > p247) ? p247 : f254;
        f255 = 2097151;
        f255 = (f255 >= `INH(p245)) ? `INH(p245) : f255;
        f255 = (f255 >= `INH(p247)) ? `INH(p247) : f255;
        f255 = (f255 > p248) ? p248 : f255;
        f256 = 2097151;
        f256 = (f256 >= `INH(p8)) ? `INH(p8) : f256;
        f256 = (f256 > p242) ? p242 : f256;
        f256 = (f256 > p246) ? p246 : f256;
        f257 = 2097151;
        f257 = (f257 > p228) ? p228 : f257;
        f257 = (f257 >= `INH(p244)) ? `INH(p244) : f257;
        f257 = (f257 >= `INH(p248)) ? `INH(p248) : f257;
        f258 = 2097151;
        f258 = (f258 > p229) ? p229 : f258;
        f258 = (f258 >= `INH(p249)) ? `INH(p249) : f258;
        f259 = 2097151;
        f259 = (f259 > p34) ? p34 : f259;
        f259 = (f259 >= `INH(p230)) ? `INH(p230) : f259;
        f260 = 2097151;
        f260 = (f260 >= `INH(p34)) ? `INH(p34) : f260;
        f260 = (f260 >= `INH(p230)) ? `INH(p230) : f260;
        f260 = (f260 > p249) ? p249 : f260;
        f261 = 2097151;
        f261 = (f261 > p9) ? p9 : f261;
        f261 = (f261 >= `INH(p229)) ? `INH(p229) : f261;
        f261 = (f261 >= `INH(p249)) ? `INH(p249) : f261;
        f262 = 2097151;
        f262 = (f262 >= `INH(p251)) ? `INH(p251) : f262;
        f262 = (f262 >= `INH(p252)) ? `INH(p252) : f262;
        f262 = (f262 > p256) ? p256 : f262;
        f263 = 2097151;
        f263 = (f263 > p250) ? p250 : f263;
        f263 = (f263 >= `INH(p256)) ? `INH(p256) : f263;
        f264 = 2097151;
        f264 = (f264 > p254) ? p254 : f264;
        f264 = (f264 >= `INH(p256)) ? `INH(p256) : f264;
        f265 = 2097151;
        f265 = (f265 >= p251/2) ? p251/2 : f265;
        f265 = (f265 >= `INH(p255)) ? `INH(p255) : f265;
        f266 = 2097151;
        f266 = (f266 >= `INH(p255)) ? `INH(p255) : f266;
        f266 = (f266 > p258) ? p258 : f266;
        f267 = 2097151;
        f267 = (f267 > p251) ? p251 : f267;
        f267 = (f267 >= `INH(p258)) ? `INH(p258) : f267;
        f267 = (f267 > p260) ? p260 : f267;
        f268 = 2097151;
        f268 = (f268 >= `INH(p258)) ? `INH(p258) : f268;
        f268 = (f268 > p261) ? p261 : f268;
        f269 = 2097151;
        f269 = (f269 > p250) ? p250 : f269;
        f269 = (f269 >= `INH(p260)) ? `INH(p260) : f269;
        f269 = (f269 >= `INH(p261)) ? `INH(p261) : f269;
        f270 = 2097151;
        f270 = (f270 > p250) ? p250 : f270;
        f270 = (f270 >= `INH(p259)) ? `INH(p259) : f270;
        f270 = (f270 >= `INH(p261)) ? `INH(p261) : f270;
        f271 = 2097151;
        f271 = (f271 >= `INH(p261)) ? `INH(p261) : f271;
        f271 = (f271 > p263) ? p263 : f271;
        f272 = 2097151;
        f272 = (f272 > p257) ? p257 : f272;
        f272 = (f272 >= `INH(p263)) ? `INH(p263) : f272;
        f273 = 2097151;
        f273 = (f273 >= `INH(p263)) ? `INH(p263) : f273;
        f273 = (f273 > p264) ? p264 : f273;
        f274 = 2097151;
        f274 = (f274 > p262) ? p262 : f274;
        f274 = (f274 >= `INH(p264)) ? `INH(p264) : f274;
        f275 = 2097151;
        f275 = (f275 > p252) ? p252 : f275;
        f275 = (f275 > p259) ? p259 : f275;
        f275 = (f275 >= `INH(p260)) ? `INH(p260) : f275;
        f275 = (f275 >= `INH(p264)) ? `INH(p264) : f275;
        f276 = 2097151;
        f276 = (f276 > p252) ? p252 : f276;
        f276 = (f276 >= `INH(p259)) ? `INH(p259) : f276;
        f276 = (f276 >= `INH(p264)) ? `INH(p264) : f276;
        f277 = 2097151;
        f277 = (f277 > p34) ? p34 : f277;
        f277 = (f277 >= `INH(p266)) ? `INH(p266) : f277;
        f278 = 2097151;
        f278 = (f278 > p265) ? p265 : f278;
        f278 = (f278 >= `INH(p267)) ? `INH(p267) : f278;
        f279 = 2097151;
        f279 = (f279 >= `INH(p34)) ? `INH(p34) : f279;
        f279 = (f279 >= `INH(p266)) ? `INH(p266) : f279;
        f279 = (f279 > p267) ? p267 : f279;
        f280 = 2097151;
        f280 = (f280 >= `INH(p265)) ? `INH(p265) : f280;
        f280 = (f280 >= `INH(p267)) ? `INH(p267) : f280;
        f280 = (f280 > p268) ? p268 : f280;
        f281 = 2097151;
        f281 = (f281 > p35) ? p35 : f281;
        f281 = (f281 >= `INH(p270)) ? `INH(p270) : f281;
        f282 = 2097151;
        f282 = (f282 > p269) ? p269 : f282;
        f282 = (f282 >= `INH(p271)) ? `INH(p271) : f282;
        f283 = 2097151;
        f283 = (f283 >= `INH(p35)) ? `INH(p35) : f283;
        f283 = (f283 >= `INH(p270)) ? `INH(p270) : f283;
        f283 = (f283 > p271) ? p271 : f283;
        f284 = 2097151;
        f284 = (f284 >= `INH(p269)) ? `INH(p269) : f284;
        f284 = (f284 >= `INH(p271)) ? `INH(p271) : f284;
        f284 = (f284 > p272) ? p272 : f284;
        f285 = 2097151;
        f285 = (f285 >= `INH(p9)) ? `INH(p9) : f285;
        f285 = (f285 > p266) ? p266 : f285;
        f285 = (f285 > p270) ? p270 : f285;
        f286 = 2097151;
        f286 = (f286 > p252) ? p252 : f286;
        f286 = (f286 >= `INH(p268)) ? `INH(p268) : f286;
        f286 = (f286 >= `INH(p272)) ? `INH(p272) : f286;
        f287 = 2097151;
        f287 = (f287 > p253) ? p253 : f287;
        f287 = (f287 >= `INH(p273)) ? `INH(p273) : f287;
        f288 = 2097151;
        f288 = (f288 > p36) ? p36 : f288;
        f288 = (f288 >= `INH(p254)) ? `INH(p254) : f288;
        f289 = 2097151;
        f289 = (f289 >= `INH(p36)) ? `INH(p36) : f289;
        f289 = (f289 >= `INH(p254)) ? `INH(p254) : f289;
        f289 = (f289 > p273) ? p273 : f289;
        f290 = 2097151;
        f290 = (f290 > p10) ? p10 : f290;
        f290 = (f290 >= `INH(p253)) ? `INH(p253) : f290;
        f290 = (f290 >= `INH(p273)) ? `INH(p273) : f290;
        f291 = 2097151;
        f291 = (f291 > p275) ? p275 : f291;
        f291 = (f291 >= `INH(p277)) ? `INH(p277) : f291;
        f292 = 2097151;
        f292 = (f292 >= `INH(p274)) ? `INH(p274) : f292;
        f292 = (f292 >= `INH(p275)) ? `INH(p275) : f292;
        f292 = (f292 >= `INH(p277)) ? `INH(p277) : f292;
        f292 = (f292 > p278) ? p278 : f292;
        f293 = 2097151;
        f293 = (f293 > p36) ? p36 : f293;
        f293 = (f293 >= `INH(p280)) ? `INH(p280) : f293;
        f294 = 2097151;
        f294 = (f294 > p279) ? p279 : f294;
        f294 = (f294 >= `INH(p281)) ? `INH(p281) : f294;
        f295 = 2097151;
        f295 = (f295 >= `INH(p36)) ? `INH(p36) : f295;
        f295 = (f295 >= `INH(p280)) ? `INH(p280) : f295;
        f295 = (f295 > p281) ? p281 : f295;
        f296 = 2097151;
        f296 = (f296 >= `INH(p279)) ? `INH(p279) : f296;
        f296 = (f296 >= `INH(p281)) ? `INH(p281) : f296;
        f296 = (f296 > p282) ? p282 : f296;
        f297 = 2097151;
        f297 = (f297 > p31) ? p31 : f297;
        f297 = (f297 >= `INH(p284)) ? `INH(p284) : f297;
        f298 = 2097151;
        f298 = (f298 > p283) ? p283 : f298;
        f298 = (f298 >= `INH(p285)) ? `INH(p285) : f298;
        f299 = 2097151;
        f299 = (f299 >= `INH(p31)) ? `INH(p31) : f299;
        f299 = (f299 >= `INH(p284)) ? `INH(p284) : f299;
        f299 = (f299 > p285) ? p285 : f299;
        f300 = 2097151;
        f300 = (f300 >= `INH(p283)) ? `INH(p283) : f300;
        f300 = (f300 >= `INH(p285)) ? `INH(p285) : f300;
        f300 = (f300 > p286) ? p286 : f300;
        f301 = 2097151;
        f301 = (f301 >= `INH(p10)) ? `INH(p10) : f301;
        f301 = (f301 > p280) ? p280 : f301;
        f301 = (f301 > p284) ? p284 : f301;
        f302 = 2097151;
        f302 = (f302 > p277) ? p277 : f302;
        f302 = (f302 >= `INH(p282)) ? `INH(p282) : f302;
        f302 = (f302 >= `INH(p286)) ? `INH(p286) : f302;
        f303 = 2097151;
        f303 = (f303 > p276) ? p276 : f303;
        f303 = (f303 >= `INH(p287)) ? `INH(p287) : f303;
        f304 = 2097151;
        f304 = (f304 > p37) ? p37 : f304;
        f304 = (f304 >= `INH(p278)) ? `INH(p278) : f304;
        f305 = 2097151;
        f305 = (f305 >= `INH(p37)) ? `INH(p37) : f305;
        f305 = (f305 >= `INH(p278)) ? `INH(p278) : f305;
        f305 = (f305 > p287) ? p287 : f305;
        f306 = 2097151;
        f306 = (f306 > p11) ? p11 : f306;
        f306 = (f306 >= `INH(p276)) ? `INH(p276) : f306;
        f306 = (f306 >= `INH(p287)) ? `INH(p287) : f306;
        f307 = 2097151;
        f307 = (f307 >= `INH(p289)) ? `INH(p289) : f307;
        f307 = (f307 >= `INH(p290)) ? `INH(p290) : f307;
        f307 = (f307 > p294) ? p294 : f307;
        f308 = 2097151;
        f308 = (f308 > p288) ? p288 : f308;
        f308 = (f308 >= `INH(p294)) ? `INH(p294) : f308;
        f309 = 2097151;
        f309 = (f309 > p292) ? p292 : f309;
        f309 = (f309 >= `INH(p294)) ? `INH(p294) : f309;
        f310 = 2097151;
        f310 = (f310 >= p289/2) ? p289/2 : f310;
        f310 = (f310 >= `INH(p293)) ? `INH(p293) : f310;
        f311 = 2097151;
        f311 = (f311 >= `INH(p293)) ? `INH(p293) : f311;
        f311 = (f311 > p296) ? p296 : f311;
        f312 = 2097151;
        f312 = (f312 > p289) ? p289 : f312;
        f312 = (f312 >= `INH(p296)) ? `INH(p296) : f312;
        f312 = (f312 > p298) ? p298 : f312;
        f313 = 2097151;
        f313 = (f313 >= `INH(p296)) ? `INH(p296) : f313;
        f313 = (f313 > p299) ? p299 : f313;
        f314 = 2097151;
        f314 = (f314 > p288) ? p288 : f314;
        f314 = (f314 >= `INH(p298)) ? `INH(p298) : f314;
        f314 = (f314 >= `INH(p299)) ? `INH(p299) : f314;
        f315 = 2097151;
        f315 = (f315 > p288) ? p288 : f315;
        f315 = (f315 >= `INH(p297)) ? `INH(p297) : f315;
        f315 = (f315 >= `INH(p299)) ? `INH(p299) : f315;
        f316 = 2097151;
        f316 = (f316 >= `INH(p299)) ? `INH(p299) : f316;
        f316 = (f316 > p301) ? p301 : f316;
        f317 = 2097151;
        f317 = (f317 > p295) ? p295 : f317;
        f317 = (f317 >= `INH(p301)) ? `INH(p301) : f317;
        f318 = 2097151;
        f318 = (f318 >= `INH(p301)) ? `INH(p301) : f318;
        f318 = (f318 > p302) ? p302 : f318;
        f319 = 2097151;
        f319 = (f319 > p300) ? p300 : f319;
        f319 = (f319 >= `INH(p302)) ? `INH(p302) : f319;
        f320 = 2097151;
        f320 = (f320 > p290) ? p290 : f320;
        f320 = (f320 > p297) ? p297 : f320;
        f320 = (f320 >= `INH(p298)) ? `INH(p298) : f320;
        f320 = (f320 >= `INH(p302)) ? `INH(p302) : f320;
        f321 = 2097151;
        f321 = (f321 > p290) ? p290 : f321;
        f321 = (f321 >= `INH(p297)) ? `INH(p297) : f321;
        f321 = (f321 >= `INH(p302)) ? `INH(p302) : f321;
        f322 = 2097151;
        f322 = (f322 > p38) ? p38 : f322;
        f322 = (f322 >= `INH(p304)) ? `INH(p304) : f322;
        f323 = 2097151;
        f323 = (f323 > p303) ? p303 : f323;
        f323 = (f323 >= `INH(p305)) ? `INH(p305) : f323;
        f324 = 2097151;
        f324 = (f324 >= `INH(p38)) ? `INH(p38) : f324;
        f324 = (f324 >= `INH(p304)) ? `INH(p304) : f324;
        f324 = (f324 > p305) ? p305 : f324;
        f325 = 2097151;
        f325 = (f325 >= `INH(p303)) ? `INH(p303) : f325;
        f325 = (f325 >= `INH(p305)) ? `INH(p305) : f325;
        f325 = (f325 > p306) ? p306 : f325;
        f326 = 2097151;
        f326 = (f326 > p39) ? p39 : f326;
        f326 = (f326 >= `INH(p308)) ? `INH(p308) : f326;
        f327 = 2097151;
        f327 = (f327 > p307) ? p307 : f327;
        f327 = (f327 >= `INH(p309)) ? `INH(p309) : f327;
        f328 = 2097151;
        f328 = (f328 >= `INH(p39)) ? `INH(p39) : f328;
        f328 = (f328 >= `INH(p308)) ? `INH(p308) : f328;
        f328 = (f328 > p309) ? p309 : f328;
        f329 = 2097151;
        f329 = (f329 >= `INH(p307)) ? `INH(p307) : f329;
        f329 = (f329 >= `INH(p309)) ? `INH(p309) : f329;
        f329 = (f329 > p310) ? p310 : f329;
        f330 = 2097151;
        f330 = (f330 >= `INH(p11)) ? `INH(p11) : f330;
        f330 = (f330 > p304) ? p304 : f330;
        f330 = (f330 > p308) ? p308 : f330;
        f331 = 2097151;
        f331 = (f331 > p290) ? p290 : f331;
        f331 = (f331 >= `INH(p306)) ? `INH(p306) : f331;
        f331 = (f331 >= `INH(p310)) ? `INH(p310) : f331;
        f332 = 2097151;
        f332 = (f332 > p291) ? p291 : f332;
        f332 = (f332 >= `INH(p311)) ? `INH(p311) : f332;
        f333 = 2097151;
        f333 = (f333 > p40) ? p40 : f333;
        f333 = (f333 >= `INH(p292)) ? `INH(p292) : f333;
        f334 = 2097151;
        f334 = (f334 >= `INH(p40)) ? `INH(p40) : f334;
        f334 = (f334 >= `INH(p292)) ? `INH(p292) : f334;
        f334 = (f334 > p311) ? p311 : f334;
        f335 = 2097151;
        f335 = (f335 > p12) ? p12 : f335;
        f335 = (f335 >= `INH(p291)) ? `INH(p291) : f335;
        f335 = (f335 >= `INH(p311)) ? `INH(p311) : f335;
        f336 = 2097151;
        f336 = (f336 > p313) ? p313 : f336;
        f336 = (f336 >= `INH(p315)) ? `INH(p315) : f336;
        f337 = 2097151;
        f337 = (f337 >= `INH(p312)) ? `INH(p312) : f337;
        f337 = (f337 >= `INH(p313)) ? `INH(p313) : f337;
        f337 = (f337 >= `INH(p315)) ? `INH(p315) : f337;
        f337 = (f337 > p316) ? p316 : f337;
        f338 = 2097151;
        f338 = (f338 > p40) ? p40 : f338;
        f338 = (f338 >= `INH(p318)) ? `INH(p318) : f338;
        f339 = 2097151;
        f339 = (f339 > p317) ? p317 : f339;
        f339 = (f339 >= `INH(p319)) ? `INH(p319) : f339;
        f340 = 2097151;
        f340 = (f340 >= `INH(p40)) ? `INH(p40) : f340;
        f340 = (f340 >= `INH(p318)) ? `INH(p318) : f340;
        f340 = (f340 > p319) ? p319 : f340;
        f341 = 2097151;
        f341 = (f341 >= `INH(p317)) ? `INH(p317) : f341;
        f341 = (f341 >= `INH(p319)) ? `INH(p319) : f341;
        f341 = (f341 > p320) ? p320 : f341;
        f342 = 2097151;
        f342 = (f342 > p37) ? p37 : f342;
        f342 = (f342 >= `INH(p322)) ? `INH(p322) : f342;
        f343 = 2097151;
        f343 = (f343 > p321) ? p321 : f343;
        f343 = (f343 >= `INH(p323)) ? `INH(p323) : f343;
        f344 = 2097151;
        f344 = (f344 >= `INH(p37)) ? `INH(p37) : f344;
        f344 = (f344 >= `INH(p322)) ? `INH(p322) : f344;
        f344 = (f344 > p323) ? p323 : f344;
        f345 = 2097151;
        f345 = (f345 >= `INH(p321)) ? `INH(p321) : f345;
        f345 = (f345 >= `INH(p323)) ? `INH(p323) : f345;
        f345 = (f345 > p324) ? p324 : f345;
        f346 = 2097151;
        f346 = (f346 >= `INH(p12)) ? `INH(p12) : f346;
        f346 = (f346 > p318) ? p318 : f346;
        f346 = (f346 > p322) ? p322 : f346;
        f347 = 2097151;
        f347 = (f347 > p315) ? p315 : f347;
        f347 = (f347 >= `INH(p320)) ? `INH(p320) : f347;
        f347 = (f347 >= `INH(p324)) ? `INH(p324) : f347;
        f348 = 2097151;
        f348 = (f348 > p314) ? p314 : f348;
        f348 = (f348 >= `INH(p325)) ? `INH(p325) : f348;
        f349 = 2097151;
        f349 = (f349 > p41) ? p41 : f349;
        f349 = (f349 >= `INH(p316)) ? `INH(p316) : f349;
        f350 = 2097151;
        f350 = (f350 >= `INH(p41)) ? `INH(p41) : f350;
        f350 = (f350 >= `INH(p316)) ? `INH(p316) : f350;
        f350 = (f350 > p325) ? p325 : f350;
        f351 = 2097151;
        f351 = (f351 > p13) ? p13 : f351;
        f351 = (f351 >= `INH(p314)) ? `INH(p314) : f351;
        f351 = (f351 >= `INH(p325)) ? `INH(p325) : f351;
        f352 = 2097151;
        f352 = (f352 > p327) ? p327 : f352;
        f352 = (f352 >= `INH(p329)) ? `INH(p329) : f352;
        f353 = 2097151;
        f353 = (f353 >= `INH(p326)) ? `INH(p326) : f353;
        f353 = (f353 >= `INH(p327)) ? `INH(p327) : f353;
        f353 = (f353 >= `INH(p329)) ? `INH(p329) : f353;
        f353 = (f353 > p330) ? p330 : f353;
        f354 = 2097151;
        f354 = (f354 > p41) ? p41 : f354;
        f354 = (f354 >= `INH(p332)) ? `INH(p332) : f354;
        f355 = 2097151;
        f355 = (f355 > p331) ? p331 : f355;
        f355 = (f355 >= `INH(p333)) ? `INH(p333) : f355;
        f356 = 2097151;
        f356 = (f356 >= `INH(p41)) ? `INH(p41) : f356;
        f356 = (f356 >= `INH(p332)) ? `INH(p332) : f356;
        f356 = (f356 > p333) ? p333 : f356;
        f357 = 2097151;
        f357 = (f357 >= `INH(p331)) ? `INH(p331) : f357;
        f357 = (f357 >= `INH(p333)) ? `INH(p333) : f357;
        f357 = (f357 > p334) ? p334 : f357;
        f358 = 2097151;
        f358 = (f358 > p42) ? p42 : f358;
        f358 = (f358 >= `INH(p336)) ? `INH(p336) : f358;
        f359 = 2097151;
        f359 = (f359 > p335) ? p335 : f359;
        f359 = (f359 >= `INH(p337)) ? `INH(p337) : f359;
        f360 = 2097151;
        f360 = (f360 >= `INH(p42)) ? `INH(p42) : f360;
        f360 = (f360 >= `INH(p336)) ? `INH(p336) : f360;
        f360 = (f360 > p337) ? p337 : f360;
        f361 = 2097151;
        f361 = (f361 >= `INH(p335)) ? `INH(p335) : f361;
        f361 = (f361 >= `INH(p337)) ? `INH(p337) : f361;
        f361 = (f361 > p338) ? p338 : f361;
        f362 = 2097151;
        f362 = (f362 >= `INH(p13)) ? `INH(p13) : f362;
        f362 = (f362 > p332) ? p332 : f362;
        f362 = (f362 > p336) ? p336 : f362;
        f363 = 2097151;
        f363 = (f363 > p329) ? p329 : f363;
        f363 = (f363 >= `INH(p334)) ? `INH(p334) : f363;
        f363 = (f363 >= `INH(p338)) ? `INH(p338) : f363;
        f364 = 2097151;
        f364 = (f364 > p328) ? p328 : f364;
        f364 = (f364 >= `INH(p339)) ? `INH(p339) : f364;
        f365 = 2097151;
        f365 = (f365 > p43) ? p43 : f365;
        f365 = (f365 >= `INH(p330)) ? `INH(p330) : f365;
        f366 = 2097151;
        f366 = (f366 >= `INH(p43)) ? `INH(p43) : f366;
        f366 = (f366 >= `INH(p330)) ? `INH(p330) : f366;
        f366 = (f366 > p339) ? p339 : f366;
        f367 = 2097151;
        f367 = (f367 > p14) ? p14 : f367;
        f367 = (f367 >= `INH(p328)) ? `INH(p328) : f367;
        f367 = (f367 >= `INH(p339)) ? `INH(p339) : f367;
        if(f14>0)
                f0 = 0;
        if(f15>0)
                f16 = 0;
        if(f17>0)
                f18 = 0;
        if(f19>0)
                f20 = 0;
        if(f21>0)
                f23 = 0;
        if(f22>0)
                f23 = 0;
        if(f24>0)
                f25 = 0;
        if(f26>0)
                f27 = 0;
        if(f26>0)
                f28 = 0;
        if(f43>0)
                f1 = 0;
        if(f44>0)
                f45 = 0;
        if(f46>0)
                f47 = 0;
        if(f48>0)
                f49 = 0;
        if(f50>0)
                f52 = 0;
        if(f51>0)
                f52 = 0;
        if(f53>0)
                f54 = 0;
        if(f55>0)
                f56 = 0;
        if(f55>0)
                f57 = 0;
        if(f72>0)
                f2 = 0;
        if(f73>0)
                f74 = 0;
        if(f75>0)
                f76 = 0;
        if(f77>0)
                f78 = 0;
        if(f79>0)
                f81 = 0;
        if(f80>0)
                f81 = 0;
        if(f82>0)
                f83 = 0;
        if(f84>0)
                f85 = 0;
        if(f84>0)
                f86 = 0;
        if(f101>0)
                f3 = 0;
        if(f102>0)
                f103 = 0;
        if(f104>0)
                f105 = 0;
        if(f106>0)
                f107 = 0;
        if(f108>0)
                f110 = 0;
        if(f109>0)
                f110 = 0;
        if(f111>0)
                f112 = 0;
        if(f113>0)
                f114 = 0;
        if(f113>0)
                f115 = 0;
        if(f130>0)
                f4 = 0;
        if(f131>0)
                f132 = 0;
        if(f133>0)
                f134 = 0;
        if(f135>0)
                f136 = 0;
        if(f137>0)
                f139 = 0;
        if(f138>0)
                f139 = 0;
        if(f140>0)
                f141 = 0;
        if(f142>0)
                f143 = 0;
        if(f142>0)
                f144 = 0;
        if(f159>0)
                f5 = 0;
        if(f160>0)
                f161 = 0;
        if(f162>0)
                f163 = 0;
        if(f164>0)
                f165 = 0;
        if(f166>0)
                f168 = 0;
        if(f167>0)
                f168 = 0;
        if(f169>0)
                f170 = 0;
        if(f171>0)
                f172 = 0;
        if(f171>0)
                f173 = 0;
        if(f188>0)
                f6 = 0;
        if(f189>0)
                f190 = 0;
        if(f191>0)
                f192 = 0;
        if(f193>0)
                f194 = 0;
        if(f195>0)
                f197 = 0;
        if(f196>0)
                f197 = 0;
        if(f198>0)
                f199 = 0;
        if(f200>0)
                f201 = 0;
        if(f200>0)
                f202 = 0;
        if(f233>0)
                f8 = 0;
        if(f234>0)
                f235 = 0;
        if(f236>0)
                f237 = 0;
        if(f238>0)
                f239 = 0;
        if(f240>0)
                f242 = 0;
        if(f241>0)
                f242 = 0;
        if(f243>0)
                f244 = 0;
        if(f245>0)
                f246 = 0;
        if(f245>0)
                f247 = 0;
        if(f262>0)
                f9 = 0;
        if(f263>0)
                f264 = 0;
        if(f265>0)
                f266 = 0;
        if(f267>0)
                f268 = 0;
        if(f269>0)
                f271 = 0;
        if(f270>0)
                f271 = 0;
        if(f272>0)
                f273 = 0;
        if(f274>0)
                f275 = 0;
        if(f274>0)
                f276 = 0;
        if(f307>0)
                f11 = 0;
        if(f308>0)
                f309 = 0;
        if(f310>0)
                f311 = 0;
        if(f312>0)
                f313 = 0;
        if(f314>0)
                f316 = 0;
        if(f315>0)
                f316 = 0;
        if(f317>0)
                f318 = 0;
        if(f319>0)
                f320 = 0;
        if(f319>0)
                f321 = 0;
        tf = (f0>0)?1:(f1>0)?2:(f2>0)?3:(f3>0)?4:(f4>0)?5:(f5>0)?6:(f6>0)?7:(f7>0)?8:(f8>0)?9:(f9>0)?10:(f10>0)?11:(f11>0)?12:(f12>0)?13:(f13>0)?14:(f14>0)?15:(f15>0)?16:(f16>0)?17:(f17>0)?18:(f18>0)?19:(f19>0)?20:(f20>0)?21:(f21>0)?22:(f22>0)?23:(f23>0)?24:(f24>0)?25:(f25>0)?26:(f26>0)?27:(f27>0)?28:(f28>0)?29:(f29>0)?30:(f30>0)?31:(f31>0)?32:(f32>0)?33:(f33>0)?34:(f34>0)?35:(f35>0)?36:(f36>0)?37:(f37>0)?38:(f38>0)?39:(f39>0)?40:(f40>0)?41:(f41>0)?42:(f42>0)?43:(f43>0)?44:(f44>0)?45:(f45>0)?46:(f46>0)?47:(f47>0)?48:(f48>0)?49:(f49>0)?50:(f50>0)?51:(f51>0)?52:(f52>0)?53:(f53>0)?54:(f54>0)?55:(f55>0)?56:(f56>0)?57:(f57>0)?58:(f58>0)?59:(f59>0)?60:(f60>0)?61:(f61>0)?62:(f62>0)?63:(f63>0)?64:(f64>0)?65:(f65>0)?66:(f66>0)?67:(f67>0)?68:(f68>0)?69:(f69>0)?70:(f70>0)?71:(f71>0)?72:(f72>0)?73:(f73>0)?74:(f74>0)?75:(f75>0)?76:(f76>0)?77:(f77>0)?78:(f78>0)?79:(f79>0)?80:(f80>0)?81:(f81>0)?82:(f82>0)?83:(f83>0)?84:(f84>0)?85:(f85>0)?86:(f86>0)?87:(f87>0)?88:(f88>0)?89:(f89>0)?90:(f90>0)?91:(f91>0)?92:(f92>0)?93:(f93>0)?94:(f94>0)?95:(f95>0)?96:(f96>0)?97:(f97>0)?98:(f98>0)?99:(f99>0)?100:(f100>0)?101:(f101>0)?102:(f102>0)?103:(f103>0)?104:(f104>0)?105:(f105>0)?106:(f106>0)?107:(f107>0)?108:(f108>0)?109:(f109>0)?110:(f110>0)?111:(f111>0)?112:(f112>0)?113:(f113>0)?114:(f114>0)?115:(f115>0)?116:(f116>0)?117:(f117>0)?118:(f118>0)?119:(f119>0)?120:(f120>0)?121:(f121>0)?122:(f122>0)?123:(f123>0)?124:(f124>0)?125:(f125>0)?126:(f126>0)?127:(f127>0)?128:(f128>0)?129:(f129>0)?130:(f130>0)?131:(f131>0)?132:(f132>0)?133:(f133>0)?134:(f134>0)?135:(f135>0)?136:(f136>0)?137:(f137>0)?138:(f138>0)?139:(f139>0)?140:(f140>0)?141:(f141>0)?142:(f142>0)?143:(f143>0)?144:(f144>0)?145:(f145>0)?146:(f146>0)?147:(f147>0)?148:(f148>0)?149:(f149>0)?150:(f150>0)?151:(f151>0)?152:(f152>0)?153:(f153>0)?154:(f154>0)?155:(f155>0)?156:(f156>0)?157:(f157>0)?158:(f158>0)?159:(f159>0)?160:(f160>0)?161:(f161>0)?162:(f162>0)?163:(f163>0)?164:(f164>0)?165:(f165>0)?166:(f166>0)?167:(f167>0)?168:(f168>0)?169:(f169>0)?170:(f170>0)?171:(f171>0)?172:(f172>0)?173:(f173>0)?174:(f174>0)?175:(f175>0)?176:(f176>0)?177:(f177>0)?178:(f178>0)?179:(f179>0)?180:(f180>0)?181:(f181>0)?182:(f182>0)?183:(f183>0)?184:(f184>0)?185:(f185>0)?186:(f186>0)?187:(f187>0)?188:(f188>0)?189:(f189>0)?190:(f190>0)?191:(f191>0)?192:(f192>0)?193:(f193>0)?194:(f194>0)?195:(f195>0)?196:(f196>0)?197:(f197>0)?198:(f198>0)?199:(f199>0)?200:(f200>0)?201:(f201>0)?202:(f202>0)?203:(f203>0)?204:(f204>0)?205:(f205>0)?206:(f206>0)?207:(f207>0)?208:(f208>0)?209:(f209>0)?210:(f210>0)?211:(f211>0)?212:(f212>0)?213:(f213>0)?214:(f214>0)?215:(f215>0)?216:(f216>0)?217:(f217>0)?218:(f218>0)?219:(f219>0)?220:(f220>0)?221:(f221>0)?222:(f222>0)?223:(f223>0)?224:(f224>0)?225:(f225>0)?226:(f226>0)?227:(f227>0)?228:(f228>0)?229:(f229>0)?230:(f230>0)?231:(f231>0)?232:(f232>0)?233:(f233>0)?234:(f234>0)?235:(f235>0)?236:(f236>0)?237:(f237>0)?238:(f238>0)?239:(f239>0)?240:(f240>0)?241:(f241>0)?242:(f242>0)?243:(f243>0)?244:(f244>0)?245:(f245>0)?246:(f246>0)?247:(f247>0)?248:(f248>0)?249:(f249>0)?250:(f250>0)?251:(f251>0)?252:(f252>0)?253:(f253>0)?254:(f254>0)?255:(f255>0)?256:(f256>0)?257:(f257>0)?258:(f258>0)?259:(f259>0)?260:(f260>0)?261:(f261>0)?262:(f262>0)?263:(f263>0)?264:(f264>0)?265:(f265>0)?266:(f266>0)?267:(f267>0)?268:(f268>0)?269:(f269>0)?270:(f270>0)?271:(f271>0)?272:(f272>0)?273:(f273>0)?274:(f274>0)?275:(f275>0)?276:(f276>0)?277:(f277>0)?278:(f278>0)?279:(f279>0)?280:(f280>0)?281:(f281>0)?282:(f282>0)?283:(f283>0)?284:(f284>0)?285:(f285>0)?286:(f286>0)?287:(f287>0)?288:(f288>0)?289:(f289>0)?290:(f290>0)?291:(f291>0)?292:(f292>0)?293:(f293>0)?294:(f294>0)?295:(f295>0)?296:(f296>0)?297:(f297>0)?298:(f298>0)?299:(f299>0)?300:(f300>0)?301:(f301>0)?302:(f302>0)?303:(f303>0)?304:(f304>0)?305:(f305>0)?306:(f306>0)?307:(f307>0)?308:(f308>0)?309:(f309>0)?310:(f310>0)?311:(f311>0)?312:(f312>0)?313:(f313>0)?314:(f314>0)?315:(f315>0)?316:(f316>0)?317:(f317>0)?318:(f318>0)?319:(f319>0)?320:(f320>0)?321:(f321>0)?322:(f322>0)?323:(f323>0)?324:(f324>0)?325:(f325>0)?326:(f326>0)?327:(f327>0)?328:(f328>0)?329:(f329>0)?330:(f330>0)?331:(f331>0)?332:(f332>0)?333:(f333>0)?334:(f334>0)?335:(f335>0)?336:(f336>0)?337:(f337>0)?338:(f338>0)?339:(f339>0)?340:(f340>0)?341:(f341>0)?342:(f342>0)?343:(f343>0)?344:(f344>0)?345:(f345>0)?346:(f346>0)?347:(f347>0)?348:(f348>0)?349:(f349>0)?350:(f350>0)?351:(f351>0)?352:(f352>0)?353:(f353>0)?354:(f354>0)?355:(f355>0)?356:(f356>0)?357:(f357>0)?358:(f358>0)?359:(f359>0)?360:(f360>0)?361:(f361>0)?362:(f362>0)?363:(f363>0)?364:(f364>0)?365:(f365>0)?366:(f366>0)?367:(f367>0)?368:0;
        case(tf)
                1: begin
                        tc = f0;
                        p49 = p49 - tc;
                        p46 = p46 + tc;
                end
                2: begin
                        tc = f1;
                        p73 = p73 - tc;
                        p70 = p70 + tc;
                end
                3: begin
                        tc = f2;
                        p97 = p97 - tc;
                        p94 = p94 + tc;
                end
                4: begin
                        tc = f3;
                        p121 = p121 - tc;
                        p118 = p118 + tc;
                end
                5: begin
                        tc = f4;
                        p145 = p145 - tc;
                        p142 = p142 + tc;
                end
                6: begin
                        tc = f5;
                        p169 = p169 - tc;
                        p166 = p166 + tc;
                end
                7: begin
                        tc = f6;
                        p193 = p193 - tc;
                        p190 = p190 + tc;
                end
                8: begin
                        tc = f7;
                        p212 = p212 - tc;
                        p214 = p214 + tc;
                end
                9: begin
                        tc = f8;
                        p231 = p231 - tc;
                        p228 = p228 + tc;
                end
                10: begin
                        tc = f9;
                        p255 = p255 - tc;
                        p252 = p252 + tc;
                end
                11: begin
                        tc = f10;
                        p274 = p274 - tc;
                        p276 = p276 + tc;
                end
                12: begin
                        tc = f11;
                        p293 = p293 - tc;
                        p290 = p290 + tc;
                end
                13: begin
                        tc = f12;
                        p312 = p312 - tc;
                        p314 = p314 + tc;
                end
                14: begin
                        tc = f13;
                        p326 = p326 - tc;
                        p328 = p328 + tc;
                end
                15: begin
                        tc = f14;
                        p50 = p50 - tc;
                        p46 = p46 + tc;
                end
                16: begin
                        tc = f15;
                        p44 = p44 - tc;
                end
                17: begin
                        tc = f16;
                        p48 = p48 - tc;
                        p50 = p50 + tc;
                end
                18: begin
                        tc = f17;
                        p45 = p45 - tc*2;
                        p51 = p51 + tc;
                end
                19: begin
                        tc = f18;
                        p52 = p52 - tc;
                        p49 = p49 + tc;
                end
                20: begin
                        tc = f19;
                        p45 = p45 - tc;
                        p54 = p54 - tc;
                        p53 = p53 + tc;
                end
                21: begin
                        tc = f20;
                        p55 = p55 - tc;
                        p52 = p52 + tc;
                end
                22: begin
                        tc = f21;
                        p44 = p44 - tc;
                        p47 = p47 + tc;
                        p56 = p56 + tc;
                end
                23: begin
                        tc = f22;
                        p44 = p44 - tc;
                        p56 = p56 + tc;
                end
                24: begin
                        tc = f23;
                        p57 = p57 - tc;
                        p55 = p55 + tc;
                end
                25: begin
                        tc = f24;
                        p51 = p51 - tc;
                        p45 = p45 + tc;
                end
                26: begin
                        tc = f25;
                        p58 = p58 - tc;
                        p57 = p57 + tc;
                end
                27: begin
                        tc = f26;
                        p56 = p56 - tc;
                        p44 = p44 + tc*2;
                end
                28: begin
                        tc = f27;
                        p46 = p46 - tc;
                        p53 = p53 - tc;
                        p54 = p54 + tc;
                        p58 = p58 + tc;
                end
                29: begin
                        tc = f28;
                        p46 = p46 - tc;
                        p58 = p58 + tc;
                end
                30: begin
                        tc = f29;
                        p15 = p15 - tc;
                        p44 = p44 + tc;
                        p59 = p59 + tc;
                end
                31: begin
                        tc = f30;
                        p59 = p59 - tc;
                        p15 = p15 + tc;
                end
                32: begin
                        tc = f31;
                        p61 = p61 - tc;
                        p60 = p60 + tc;
                end
                33: begin
                        tc = f32;
                        p62 = p62 - tc;
                        p61 = p61 + tc;
                end
                34: begin
                        tc = f33;
                        p16 = p16 - tc;
                        p45 = p45 + tc;
                        p63 = p63 + tc;
                end
                35: begin
                        tc = f34;
                        p63 = p63 - tc;
                        p16 = p16 + tc;
                end
                36: begin
                        tc = f35;
                        p65 = p65 - tc;
                        p64 = p64 + tc;
                end
                37: begin
                        tc = f36;
                        p66 = p66 - tc;
                        p65 = p65 + tc;
                end
                38: begin
                        tc = f37;
                        p60 = p60 - tc;
                        p64 = p64 - tc;
                        p0 = p0 + tc;
                end
                39: begin
                        tc = f38;
                        p46 = p46 - tc;
                        p62 = p62 + tc;
                        p66 = p66 + tc;
                end
                40: begin
                        tc = f39;
                        p47 = p47 - tc;
                        p17 = p17 + tc;
                end
                41: begin
                        tc = f40;
                        p17 = p17 - tc;
                end
                42: begin
                        tc = f41;
                        p67 = p67 - tc;
                        p48 = p48 + tc;
                end
                43: begin
                        tc = f42;
                        p1 = p1 - tc;
                        p67 = p67 + tc;
                end
                44: begin
                        tc = f43;
                        p74 = p74 - tc;
                        p70 = p70 + tc;
                end
                45: begin
                        tc = f44;
                        p68 = p68 - tc;
                end
                46: begin
                        tc = f45;
                        p72 = p72 - tc;
                        p74 = p74 + tc;
                end
                47: begin
                        tc = f46;
                        p69 = p69 - tc*2;
                        p75 = p75 + tc;
                end
                48: begin
                        tc = f47;
                        p76 = p76 - tc;
                        p73 = p73 + tc;
                end
                49: begin
                        tc = f48;
                        p69 = p69 - tc;
                        p78 = p78 - tc;
                        p77 = p77 + tc;
                end
                50: begin
                        tc = f49;
                        p79 = p79 - tc;
                        p76 = p76 + tc;
                end
                51: begin
                        tc = f50;
                        p68 = p68 - tc;
                        p71 = p71 + tc;
                        p80 = p80 + tc;
                end
                52: begin
                        tc = f51;
                        p68 = p68 - tc;
                        p80 = p80 + tc;
                end
                53: begin
                        tc = f52;
                        p81 = p81 - tc;
                        p79 = p79 + tc;
                end
                54: begin
                        tc = f53;
                        p75 = p75 - tc;
                        p69 = p69 + tc;
                end
                55: begin
                        tc = f54;
                        p82 = p82 - tc;
                        p81 = p81 + tc;
                end
                56: begin
                        tc = f55;
                        p80 = p80 - tc;
                        p68 = p68 + tc*2;
                end
                57: begin
                        tc = f56;
                        p70 = p70 - tc;
                        p77 = p77 - tc;
                        p78 = p78 + tc;
                        p82 = p82 + tc;
                end
                58: begin
                        tc = f57;
                        p70 = p70 - tc;
                        p82 = p82 + tc;
                end
                59: begin
                        tc = f58;
                        p17 = p17 - tc;
                        p68 = p68 + tc;
                        p83 = p83 + tc;
                end
                60: begin
                        tc = f59;
                        p83 = p83 - tc;
                        p17 = p17 + tc;
                end
                61: begin
                        tc = f60;
                        p85 = p85 - tc;
                        p84 = p84 + tc;
                end
                62: begin
                        tc = f61;
                        p86 = p86 - tc;
                        p85 = p85 + tc;
                end
                63: begin
                        tc = f62;
                        p18 = p18 - tc;
                        p69 = p69 + tc;
                        p87 = p87 + tc;
                end
                64: begin
                        tc = f63;
                        p87 = p87 - tc;
                        p18 = p18 + tc;
                end
                65: begin
                        tc = f64;
                        p89 = p89 - tc;
                        p88 = p88 + tc;
                end
                66: begin
                        tc = f65;
                        p90 = p90 - tc;
                        p89 = p89 + tc;
                end
                67: begin
                        tc = f66;
                        p84 = p84 - tc;
                        p88 = p88 - tc;
                        p1 = p1 + tc;
                end
                68: begin
                        tc = f67;
                        p70 = p70 - tc;
                        p86 = p86 + tc;
                        p90 = p90 + tc;
                end
                69: begin
                        tc = f68;
                        p71 = p71 - tc;
                        p19 = p19 + tc;
                end
                70: begin
                        tc = f69;
                        p19 = p19 - tc;
                end
                71: begin
                        tc = f70;
                        p91 = p91 - tc;
                        p72 = p72 + tc;
                end
                72: begin
                        tc = f71;
                        p2 = p2 - tc;
                        p91 = p91 + tc;
                end
                73: begin
                        tc = f72;
                        p98 = p98 - tc;
                        p94 = p94 + tc;
                end
                74: begin
                        tc = f73;
                        p92 = p92 - tc;
                end
                75: begin
                        tc = f74;
                        p96 = p96 - tc;
                        p98 = p98 + tc;
                end
                76: begin
                        tc = f75;
                        p93 = p93 - tc*2;
                        p99 = p99 + tc;
                end
                77: begin
                        tc = f76;
                        p100 = p100 - tc;
                        p97 = p97 + tc;
                end
                78: begin
                        tc = f77;
                        p93 = p93 - tc;
                        p102 = p102 - tc;
                        p101 = p101 + tc;
                end
                79: begin
                        tc = f78;
                        p103 = p103 - tc;
                        p100 = p100 + tc;
                end
                80: begin
                        tc = f79;
                        p92 = p92 - tc;
                        p95 = p95 + tc;
                        p104 = p104 + tc;
                end
                81: begin
                        tc = f80;
                        p92 = p92 - tc;
                        p104 = p104 + tc;
                end
                82: begin
                        tc = f81;
                        p105 = p105 - tc;
                        p103 = p103 + tc;
                end
                83: begin
                        tc = f82;
                        p99 = p99 - tc;
                        p93 = p93 + tc;
                end
                84: begin
                        tc = f83;
                        p106 = p106 - tc;
                        p105 = p105 + tc;
                end
                85: begin
                        tc = f84;
                        p104 = p104 - tc;
                        p92 = p92 + tc*2;
                end
                86: begin
                        tc = f85;
                        p94 = p94 - tc;
                        p101 = p101 - tc;
                        p102 = p102 + tc;
                        p106 = p106 + tc;
                end
                87: begin
                        tc = f86;
                        p94 = p94 - tc;
                        p106 = p106 + tc;
                end
                88: begin
                        tc = f87;
                        p19 = p19 - tc;
                        p92 = p92 + tc;
                        p107 = p107 + tc;
                end
                89: begin
                        tc = f88;
                        p107 = p107 - tc;
                        p19 = p19 + tc;
                end
                90: begin
                        tc = f89;
                        p109 = p109 - tc;
                        p108 = p108 + tc;
                end
                91: begin
                        tc = f90;
                        p110 = p110 - tc;
                        p109 = p109 + tc;
                end
                92: begin
                        tc = f91;
                        p20 = p20 - tc;
                        p93 = p93 + tc;
                        p111 = p111 + tc;
                end
                93: begin
                        tc = f92;
                        p111 = p111 - tc;
                        p20 = p20 + tc;
                end
                94: begin
                        tc = f93;
                        p113 = p113 - tc;
                        p112 = p112 + tc;
                end
                95: begin
                        tc = f94;
                        p114 = p114 - tc;
                        p113 = p113 + tc;
                end
                96: begin
                        tc = f95;
                        p108 = p108 - tc;
                        p112 = p112 - tc;
                        p2 = p2 + tc;
                end
                97: begin
                        tc = f96;
                        p94 = p94 - tc;
                        p110 = p110 + tc;
                        p114 = p114 + tc;
                end
                98: begin
                        tc = f97;
                        p95 = p95 - tc;
                        p21 = p21 + tc;
                end
                99: begin
                        tc = f98;
                        p21 = p21 - tc;
                end
                100: begin
                        tc = f99;
                        p115 = p115 - tc;
                        p96 = p96 + tc;
                end
                101: begin
                        tc = f100;
                        p3 = p3 - tc;
                        p115 = p115 + tc;
                end
                102: begin
                        tc = f101;
                        p122 = p122 - tc;
                        p118 = p118 + tc;
                end
                103: begin
                        tc = f102;
                        p116 = p116 - tc;
                end
                104: begin
                        tc = f103;
                        p120 = p120 - tc;
                        p122 = p122 + tc;
                end
                105: begin
                        tc = f104;
                        p117 = p117 - tc*2;
                        p123 = p123 + tc;
                end
                106: begin
                        tc = f105;
                        p124 = p124 - tc;
                        p121 = p121 + tc;
                end
                107: begin
                        tc = f106;
                        p117 = p117 - tc;
                        p126 = p126 - tc;
                        p125 = p125 + tc;
                end
                108: begin
                        tc = f107;
                        p127 = p127 - tc;
                        p124 = p124 + tc;
                end
                109: begin
                        tc = f108;
                        p116 = p116 - tc;
                        p119 = p119 + tc;
                        p128 = p128 + tc;
                end
                110: begin
                        tc = f109;
                        p116 = p116 - tc;
                        p128 = p128 + tc;
                end
                111: begin
                        tc = f110;
                        p129 = p129 - tc;
                        p127 = p127 + tc;
                end
                112: begin
                        tc = f111;
                        p123 = p123 - tc;
                        p117 = p117 + tc;
                end
                113: begin
                        tc = f112;
                        p130 = p130 - tc;
                        p129 = p129 + tc;
                end
                114: begin
                        tc = f113;
                        p128 = p128 - tc;
                        p116 = p116 + tc*2;
                end
                115: begin
                        tc = f114;
                        p118 = p118 - tc;
                        p125 = p125 - tc;
                        p126 = p126 + tc;
                        p130 = p130 + tc;
                end
                116: begin
                        tc = f115;
                        p118 = p118 - tc;
                        p130 = p130 + tc;
                end
                117: begin
                        tc = f116;
                        p21 = p21 - tc;
                        p116 = p116 + tc;
                        p131 = p131 + tc;
                end
                118: begin
                        tc = f117;
                        p131 = p131 - tc;
                        p21 = p21 + tc;
                end
                119: begin
                        tc = f118;
                        p133 = p133 - tc;
                        p132 = p132 + tc;
                end
                120: begin
                        tc = f119;
                        p134 = p134 - tc;
                        p133 = p133 + tc;
                end
                121: begin
                        tc = f120;
                        p22 = p22 - tc;
                        p117 = p117 + tc;
                        p135 = p135 + tc;
                end
                122: begin
                        tc = f121;
                        p135 = p135 - tc;
                        p22 = p22 + tc;
                end
                123: begin
                        tc = f122;
                        p137 = p137 - tc;
                        p136 = p136 + tc;
                end
                124: begin
                        tc = f123;
                        p138 = p138 - tc;
                        p137 = p137 + tc;
                end
                125: begin
                        tc = f124;
                        p132 = p132 - tc;
                        p136 = p136 - tc;
                        p3 = p3 + tc;
                end
                126: begin
                        tc = f125;
                        p118 = p118 - tc;
                        p134 = p134 + tc;
                        p138 = p138 + tc;
                end
                127: begin
                        tc = f126;
                        p119 = p119 - tc;
                        p23 = p23 + tc;
                end
                128: begin
                        tc = f127;
                        p23 = p23 - tc;
                end
                129: begin
                        tc = f128;
                        p139 = p139 - tc;
                        p120 = p120 + tc;
                end
                130: begin
                        tc = f129;
                        p4 = p4 - tc;
                        p139 = p139 + tc;
                end
                131: begin
                        tc = f130;
                        p146 = p146 - tc;
                        p142 = p142 + tc;
                end
                132: begin
                        tc = f131;
                        p140 = p140 - tc;
                end
                133: begin
                        tc = f132;
                        p144 = p144 - tc;
                        p146 = p146 + tc;
                end
                134: begin
                        tc = f133;
                        p141 = p141 - tc*2;
                        p147 = p147 + tc;
                end
                135: begin
                        tc = f134;
                        p148 = p148 - tc;
                        p145 = p145 + tc;
                end
                136: begin
                        tc = f135;
                        p141 = p141 - tc;
                        p150 = p150 - tc;
                        p149 = p149 + tc;
                end
                137: begin
                        tc = f136;
                        p151 = p151 - tc;
                        p148 = p148 + tc;
                end
                138: begin
                        tc = f137;
                        p140 = p140 - tc;
                        p143 = p143 + tc;
                        p152 = p152 + tc;
                end
                139: begin
                        tc = f138;
                        p140 = p140 - tc;
                        p152 = p152 + tc;
                end
                140: begin
                        tc = f139;
                        p153 = p153 - tc;
                        p151 = p151 + tc;
                end
                141: begin
                        tc = f140;
                        p147 = p147 - tc;
                        p141 = p141 + tc;
                end
                142: begin
                        tc = f141;
                        p154 = p154 - tc;
                        p153 = p153 + tc;
                end
                143: begin
                        tc = f142;
                        p152 = p152 - tc;
                        p140 = p140 + tc*2;
                end
                144: begin
                        tc = f143;
                        p142 = p142 - tc;
                        p149 = p149 - tc;
                        p150 = p150 + tc;
                        p154 = p154 + tc;
                end
                145: begin
                        tc = f144;
                        p142 = p142 - tc;
                        p154 = p154 + tc;
                end
                146: begin
                        tc = f145;
                        p24 = p24 - tc;
                        p140 = p140 + tc;
                        p155 = p155 + tc;
                end
                147: begin
                        tc = f146;
                        p155 = p155 - tc;
                        p24 = p24 + tc;
                end
                148: begin
                        tc = f147;
                        p157 = p157 - tc;
                        p156 = p156 + tc;
                end
                149: begin
                        tc = f148;
                        p158 = p158 - tc;
                        p157 = p157 + tc;
                end
                150: begin
                        tc = f149;
                        p25 = p25 - tc;
                        p141 = p141 + tc;
                        p159 = p159 + tc;
                end
                151: begin
                        tc = f150;
                        p159 = p159 - tc;
                        p25 = p25 + tc;
                end
                152: begin
                        tc = f151;
                        p161 = p161 - tc;
                        p160 = p160 + tc;
                end
                153: begin
                        tc = f152;
                        p162 = p162 - tc;
                        p161 = p161 + tc;
                end
                154: begin
                        tc = f153;
                        p156 = p156 - tc;
                        p160 = p160 - tc;
                        p4 = p4 + tc;
                end
                155: begin
                        tc = f154;
                        p142 = p142 - tc;
                        p158 = p158 + tc;
                        p162 = p162 + tc;
                end
                156: begin
                        tc = f155;
                        p143 = p143 - tc;
                        p26 = p26 + tc;
                end
                157: begin
                        tc = f156;
                        p26 = p26 - tc;
                end
                158: begin
                        tc = f157;
                        p163 = p163 - tc;
                        p144 = p144 + tc;
                end
                159: begin
                        tc = f158;
                        p5 = p5 - tc;
                        p163 = p163 + tc;
                end
                160: begin
                        tc = f159;
                        p170 = p170 - tc;
                        p166 = p166 + tc;
                end
                161: begin
                        tc = f160;
                        p164 = p164 - tc;
                end
                162: begin
                        tc = f161;
                        p168 = p168 - tc;
                        p170 = p170 + tc;
                end
                163: begin
                        tc = f162;
                        p165 = p165 - tc*2;
                        p171 = p171 + tc;
                end
                164: begin
                        tc = f163;
                        p172 = p172 - tc;
                        p169 = p169 + tc;
                end
                165: begin
                        tc = f164;
                        p165 = p165 - tc;
                        p174 = p174 - tc;
                        p173 = p173 + tc;
                end
                166: begin
                        tc = f165;
                        p175 = p175 - tc;
                        p172 = p172 + tc;
                end
                167: begin
                        tc = f166;
                        p164 = p164 - tc;
                        p167 = p167 + tc;
                        p176 = p176 + tc;
                end
                168: begin
                        tc = f167;
                        p164 = p164 - tc;
                        p176 = p176 + tc;
                end
                169: begin
                        tc = f168;
                        p177 = p177 - tc;
                        p175 = p175 + tc;
                end
                170: begin
                        tc = f169;
                        p171 = p171 - tc;
                        p165 = p165 + tc;
                end
                171: begin
                        tc = f170;
                        p178 = p178 - tc;
                        p177 = p177 + tc;
                end
                172: begin
                        tc = f171;
                        p176 = p176 - tc;
                        p164 = p164 + tc*2;
                end
                173: begin
                        tc = f172;
                        p166 = p166 - tc;
                        p173 = p173 - tc;
                        p174 = p174 + tc;
                        p178 = p178 + tc;
                end
                174: begin
                        tc = f173;
                        p166 = p166 - tc;
                        p178 = p178 + tc;
                end
                175: begin
                        tc = f174;
                        p26 = p26 - tc;
                        p164 = p164 + tc;
                        p179 = p179 + tc;
                end
                176: begin
                        tc = f175;
                        p179 = p179 - tc;
                        p26 = p26 + tc;
                end
                177: begin
                        tc = f176;
                        p181 = p181 - tc;
                        p180 = p180 + tc;
                end
                178: begin
                        tc = f177;
                        p182 = p182 - tc;
                        p181 = p181 + tc;
                end
                179: begin
                        tc = f178;
                        p27 = p27 - tc;
                        p165 = p165 + tc;
                        p183 = p183 + tc;
                end
                180: begin
                        tc = f179;
                        p183 = p183 - tc;
                        p27 = p27 + tc;
                end
                181: begin
                        tc = f180;
                        p185 = p185 - tc;
                        p184 = p184 + tc;
                end
                182: begin
                        tc = f181;
                        p186 = p186 - tc;
                        p185 = p185 + tc;
                end
                183: begin
                        tc = f182;
                        p180 = p180 - tc;
                        p184 = p184 - tc;
                        p5 = p5 + tc;
                end
                184: begin
                        tc = f183;
                        p166 = p166 - tc;
                        p182 = p182 + tc;
                        p186 = p186 + tc;
                end
                185: begin
                        tc = f184;
                        p167 = p167 - tc;
                        p28 = p28 + tc;
                end
                186: begin
                        tc = f185;
                        p28 = p28 - tc;
                end
                187: begin
                        tc = f186;
                        p187 = p187 - tc;
                        p168 = p168 + tc;
                end
                188: begin
                        tc = f187;
                        p6 = p6 - tc;
                        p187 = p187 + tc;
                end
                189: begin
                        tc = f188;
                        p194 = p194 - tc;
                        p190 = p190 + tc;
                end
                190: begin
                        tc = f189;
                        p188 = p188 - tc;
                end
                191: begin
                        tc = f190;
                        p192 = p192 - tc;
                        p194 = p194 + tc;
                end
                192: begin
                        tc = f191;
                        p189 = p189 - tc*2;
                        p195 = p195 + tc;
                end
                193: begin
                        tc = f192;
                        p196 = p196 - tc;
                        p193 = p193 + tc;
                end
                194: begin
                        tc = f193;
                        p189 = p189 - tc;
                        p198 = p198 - tc;
                        p197 = p197 + tc;
                end
                195: begin
                        tc = f194;
                        p199 = p199 - tc;
                        p196 = p196 + tc;
                end
                196: begin
                        tc = f195;
                        p188 = p188 - tc;
                        p191 = p191 + tc;
                        p200 = p200 + tc;
                end
                197: begin
                        tc = f196;
                        p188 = p188 - tc;
                        p200 = p200 + tc;
                end
                198: begin
                        tc = f197;
                        p201 = p201 - tc;
                        p199 = p199 + tc;
                end
                199: begin
                        tc = f198;
                        p195 = p195 - tc;
                        p189 = p189 + tc;
                end
                200: begin
                        tc = f199;
                        p202 = p202 - tc;
                        p201 = p201 + tc;
                end
                201: begin
                        tc = f200;
                        p200 = p200 - tc;
                        p188 = p188 + tc*2;
                end
                202: begin
                        tc = f201;
                        p190 = p190 - tc;
                        p197 = p197 - tc;
                        p198 = p198 + tc;
                        p202 = p202 + tc;
                end
                203: begin
                        tc = f202;
                        p190 = p190 - tc;
                        p202 = p202 + tc;
                end
                204: begin
                        tc = f203;
                        p28 = p28 - tc;
                        p188 = p188 + tc;
                        p203 = p203 + tc;
                end
                205: begin
                        tc = f204;
                        p203 = p203 - tc;
                        p28 = p28 + tc;
                end
                206: begin
                        tc = f205;
                        p205 = p205 - tc;
                        p204 = p204 + tc;
                end
                207: begin
                        tc = f206;
                        p206 = p206 - tc;
                        p205 = p205 + tc;
                end
                208: begin
                        tc = f207;
                        p29 = p29 - tc;
                        p189 = p189 + tc;
                        p207 = p207 + tc;
                end
                209: begin
                        tc = f208;
                        p207 = p207 - tc;
                        p29 = p29 + tc;
                end
                210: begin
                        tc = f209;
                        p209 = p209 - tc;
                        p208 = p208 + tc;
                end
                211: begin
                        tc = f210;
                        p210 = p210 - tc;
                        p209 = p209 + tc;
                end
                212: begin
                        tc = f211;
                        p204 = p204 - tc;
                        p208 = p208 - tc;
                        p6 = p6 + tc;
                end
                213: begin
                        tc = f212;
                        p190 = p190 - tc;
                        p206 = p206 + tc;
                        p210 = p210 + tc;
                end
                214: begin
                        tc = f213;
                        p191 = p191 - tc;
                        p30 = p30 + tc;
                end
                215: begin
                        tc = f214;
                        p30 = p30 - tc;
                end
                216: begin
                        tc = f215;
                        p211 = p211 - tc;
                        p192 = p192 + tc;
                end
                217: begin
                        tc = f216;
                        p7 = p7 - tc;
                        p211 = p211 + tc;
                end
                218: begin
                        tc = f217;
                        p213 = p213 - tc;
                        p214 = p214 + tc;
                end
                219: begin
                        tc = f218;
                        p216 = p216 - tc;
                        p215 = p215 + tc;
                end
                220: begin
                        tc = f219;
                        p23 = p23 - tc;
                        p212 = p212 + tc;
                        p217 = p217 + tc;
                end
                221: begin
                        tc = f220;
                        p217 = p217 - tc;
                        p23 = p23 + tc;
                end
                222: begin
                        tc = f221;
                        p219 = p219 - tc;
                        p218 = p218 + tc;
                end
                223: begin
                        tc = f222;
                        p220 = p220 - tc;
                        p219 = p219 + tc;
                end
                224: begin
                        tc = f223;
                        p30 = p30 - tc;
                        p213 = p213 + tc;
                        p221 = p221 + tc;
                end
                225: begin
                        tc = f224;
                        p221 = p221 - tc;
                        p30 = p30 + tc;
                end
                226: begin
                        tc = f225;
                        p223 = p223 - tc;
                        p222 = p222 + tc;
                end
                227: begin
                        tc = f226;
                        p224 = p224 - tc;
                        p223 = p223 + tc;
                end
                228: begin
                        tc = f227;
                        p218 = p218 - tc;
                        p222 = p222 - tc;
                        p7 = p7 + tc;
                end
                229: begin
                        tc = f228;
                        p215 = p215 - tc;
                        p220 = p220 + tc;
                        p224 = p224 + tc;
                end
                230: begin
                        tc = f229;
                        p214 = p214 - tc;
                        p31 = p31 + tc;
                end
                231: begin
                        tc = f230;
                        p31 = p31 - tc;
                end
                232: begin
                        tc = f231;
                        p225 = p225 - tc;
                        p216 = p216 + tc;
                end
                233: begin
                        tc = f232;
                        p8 = p8 - tc;
                        p225 = p225 + tc;
                end
                234: begin
                        tc = f233;
                        p232 = p232 - tc;
                        p228 = p228 + tc;
                end
                235: begin
                        tc = f234;
                        p226 = p226 - tc;
                end
                236: begin
                        tc = f235;
                        p230 = p230 - tc;
                        p232 = p232 + tc;
                end
                237: begin
                        tc = f236;
                        p227 = p227 - tc*2;
                        p233 = p233 + tc;
                end
                238: begin
                        tc = f237;
                        p234 = p234 - tc;
                        p231 = p231 + tc;
                end
                239: begin
                        tc = f238;
                        p227 = p227 - tc;
                        p236 = p236 - tc;
                        p235 = p235 + tc;
                end
                240: begin
                        tc = f239;
                        p237 = p237 - tc;
                        p234 = p234 + tc;
                end
                241: begin
                        tc = f240;
                        p226 = p226 - tc;
                        p229 = p229 + tc;
                        p238 = p238 + tc;
                end
                242: begin
                        tc = f241;
                        p226 = p226 - tc;
                        p238 = p238 + tc;
                end
                243: begin
                        tc = f242;
                        p239 = p239 - tc;
                        p237 = p237 + tc;
                end
                244: begin
                        tc = f243;
                        p233 = p233 - tc;
                        p227 = p227 + tc;
                end
                245: begin
                        tc = f244;
                        p240 = p240 - tc;
                        p239 = p239 + tc;
                end
                246: begin
                        tc = f245;
                        p238 = p238 - tc;
                        p226 = p226 + tc*2;
                end
                247: begin
                        tc = f246;
                        p228 = p228 - tc;
                        p235 = p235 - tc;
                        p236 = p236 + tc;
                        p240 = p240 + tc;
                end
                248: begin
                        tc = f247;
                        p228 = p228 - tc;
                        p240 = p240 + tc;
                end
                249: begin
                        tc = f248;
                        p32 = p32 - tc;
                        p226 = p226 + tc;
                        p241 = p241 + tc;
                end
                250: begin
                        tc = f249;
                        p241 = p241 - tc;
                        p32 = p32 + tc;
                end
                251: begin
                        tc = f250;
                        p243 = p243 - tc;
                        p242 = p242 + tc;
                end
                252: begin
                        tc = f251;
                        p244 = p244 - tc;
                        p243 = p243 + tc;
                end
                253: begin
                        tc = f252;
                        p33 = p33 - tc;
                        p227 = p227 + tc;
                        p245 = p245 + tc;
                end
                254: begin
                        tc = f253;
                        p245 = p245 - tc;
                        p33 = p33 + tc;
                end
                255: begin
                        tc = f254;
                        p247 = p247 - tc;
                        p246 = p246 + tc;
                end
                256: begin
                        tc = f255;
                        p248 = p248 - tc;
                        p247 = p247 + tc;
                end
                257: begin
                        tc = f256;
                        p242 = p242 - tc;
                        p246 = p246 - tc;
                        p8 = p8 + tc;
                end
                258: begin
                        tc = f257;
                        p228 = p228 - tc;
                        p244 = p244 + tc;
                        p248 = p248 + tc;
                end
                259: begin
                        tc = f258;
                        p229 = p229 - tc;
                        p34 = p34 + tc;
                end
                260: begin
                        tc = f259;
                        p34 = p34 - tc;
                end
                261: begin
                        tc = f260;
                        p249 = p249 - tc;
                        p230 = p230 + tc;
                end
                262: begin
                        tc = f261;
                        p9 = p9 - tc;
                        p249 = p249 + tc;
                end
                263: begin
                        tc = f262;
                        p256 = p256 - tc;
                        p252 = p252 + tc;
                end
                264: begin
                        tc = f263;
                        p250 = p250 - tc;
                end
                265: begin
                        tc = f264;
                        p254 = p254 - tc;
                        p256 = p256 + tc;
                end
                266: begin
                        tc = f265;
                        p251 = p251 - tc*2;
                        p257 = p257 + tc;
                end
                267: begin
                        tc = f266;
                        p258 = p258 - tc;
                        p255 = p255 + tc;
                end
                268: begin
                        tc = f267;
                        p251 = p251 - tc;
                        p260 = p260 - tc;
                        p259 = p259 + tc;
                end
                269: begin
                        tc = f268;
                        p261 = p261 - tc;
                        p258 = p258 + tc;
                end
                270: begin
                        tc = f269;
                        p250 = p250 - tc;
                        p253 = p253 + tc;
                        p262 = p262 + tc;
                end
                271: begin
                        tc = f270;
                        p250 = p250 - tc;
                        p262 = p262 + tc;
                end
                272: begin
                        tc = f271;
                        p263 = p263 - tc;
                        p261 = p261 + tc;
                end
                273: begin
                        tc = f272;
                        p257 = p257 - tc;
                        p251 = p251 + tc;
                end
                274: begin
                        tc = f273;
                        p264 = p264 - tc;
                        p263 = p263 + tc;
                end
                275: begin
                        tc = f274;
                        p262 = p262 - tc;
                        p250 = p250 + tc*2;
                end
                276: begin
                        tc = f275;
                        p252 = p252 - tc;
                        p259 = p259 - tc;
                        p260 = p260 + tc;
                        p264 = p264 + tc;
                end
                277: begin
                        tc = f276;
                        p252 = p252 - tc;
                        p264 = p264 + tc;
                end
                278: begin
                        tc = f277;
                        p34 = p34 - tc;
                        p250 = p250 + tc;
                        p265 = p265 + tc;
                end
                279: begin
                        tc = f278;
                        p265 = p265 - tc;
                        p34 = p34 + tc;
                end
                280: begin
                        tc = f279;
                        p267 = p267 - tc;
                        p266 = p266 + tc;
                end
                281: begin
                        tc = f280;
                        p268 = p268 - tc;
                        p267 = p267 + tc;
                end
                282: begin
                        tc = f281;
                        p35 = p35 - tc;
                        p251 = p251 + tc;
                        p269 = p269 + tc;
                end
                283: begin
                        tc = f282;
                        p269 = p269 - tc;
                        p35 = p35 + tc;
                end
                284: begin
                        tc = f283;
                        p271 = p271 - tc;
                        p270 = p270 + tc;
                end
                285: begin
                        tc = f284;
                        p272 = p272 - tc;
                        p271 = p271 + tc;
                end
                286: begin
                        tc = f285;
                        p266 = p266 - tc;
                        p270 = p270 - tc;
                        p9 = p9 + tc;
                end
                287: begin
                        tc = f286;
                        p252 = p252 - tc;
                        p268 = p268 + tc;
                        p272 = p272 + tc;
                end
                288: begin
                        tc = f287;
                        p253 = p253 - tc;
                        p36 = p36 + tc;
                end
                289: begin
                        tc = f288;
                        p36 = p36 - tc;
                end
                290: begin
                        tc = f289;
                        p273 = p273 - tc;
                        p254 = p254 + tc;
                end
                291: begin
                        tc = f290;
                        p10 = p10 - tc;
                        p273 = p273 + tc;
                end
                292: begin
                        tc = f291;
                        p275 = p275 - tc;
                        p276 = p276 + tc;
                end
                293: begin
                        tc = f292;
                        p278 = p278 - tc;
                        p277 = p277 + tc;
                end
                294: begin
                        tc = f293;
                        p36 = p36 - tc;
                        p274 = p274 + tc;
                        p279 = p279 + tc;
                end
                295: begin
                        tc = f294;
                        p279 = p279 - tc;
                        p36 = p36 + tc;
                end
                296: begin
                        tc = f295;
                        p281 = p281 - tc;
                        p280 = p280 + tc;
                end
                297: begin
                        tc = f296;
                        p282 = p282 - tc;
                        p281 = p281 + tc;
                end
                298: begin
                        tc = f297;
                        p31 = p31 - tc;
                        p275 = p275 + tc;
                        p283 = p283 + tc;
                end
                299: begin
                        tc = f298;
                        p283 = p283 - tc;
                        p31 = p31 + tc;
                end
                300: begin
                        tc = f299;
                        p285 = p285 - tc;
                        p284 = p284 + tc;
                end
                301: begin
                        tc = f300;
                        p286 = p286 - tc;
                        p285 = p285 + tc;
                end
                302: begin
                        tc = f301;
                        p280 = p280 - tc;
                        p284 = p284 - tc;
                        p10 = p10 + tc;
                end
                303: begin
                        tc = f302;
                        p277 = p277 - tc;
                        p282 = p282 + tc;
                        p286 = p286 + tc;
                end
                304: begin
                        tc = f303;
                        p276 = p276 - tc;
                        p37 = p37 + tc;
                end
                305: begin
                        tc = f304;
                        p37 = p37 - tc;
                end
                306: begin
                        tc = f305;
                        p287 = p287 - tc;
                        p278 = p278 + tc;
                end
                307: begin
                        tc = f306;
                        p11 = p11 - tc;
                        p287 = p287 + tc;
                end
                308: begin
                        tc = f307;
                        p294 = p294 - tc;
                        p290 = p290 + tc;
                end
                309: begin
                        tc = f308;
                        p288 = p288 - tc;
                end
                310: begin
                        tc = f309;
                        p292 = p292 - tc;
                        p294 = p294 + tc;
                end
                311: begin
                        tc = f310;
                        p289 = p289 - tc*2;
                        p295 = p295 + tc;
                end
                312: begin
                        tc = f311;
                        p296 = p296 - tc;
                        p293 = p293 + tc;
                end
                313: begin
                        tc = f312;
                        p289 = p289 - tc;
                        p298 = p298 - tc;
                        p297 = p297 + tc;
                end
                314: begin
                        tc = f313;
                        p299 = p299 - tc;
                        p296 = p296 + tc;
                end
                315: begin
                        tc = f314;
                        p288 = p288 - tc;
                        p291 = p291 + tc;
                        p300 = p300 + tc;
                end
                316: begin
                        tc = f315;
                        p288 = p288 - tc;
                        p300 = p300 + tc;
                end
                317: begin
                        tc = f316;
                        p301 = p301 - tc;
                        p299 = p299 + tc;
                end
                318: begin
                        tc = f317;
                        p295 = p295 - tc;
                        p289 = p289 + tc;
                end
                319: begin
                        tc = f318;
                        p302 = p302 - tc;
                        p301 = p301 + tc;
                end
                320: begin
                        tc = f319;
                        p300 = p300 - tc;
                        p288 = p288 + tc*2;
                end
                321: begin
                        tc = f320;
                        p290 = p290 - tc;
                        p297 = p297 - tc;
                        p298 = p298 + tc;
                        p302 = p302 + tc;
                end
                322: begin
                        tc = f321;
                        p290 = p290 - tc;
                        p302 = p302 + tc;
                end
                323: begin
                        tc = f322;
                        p38 = p38 - tc;
                        p288 = p288 + tc;
                        p303 = p303 + tc;
                end
                324: begin
                        tc = f323;
                        p303 = p303 - tc;
                        p38 = p38 + tc;
                end
                325: begin
                        tc = f324;
                        p305 = p305 - tc;
                        p304 = p304 + tc;
                end
                326: begin
                        tc = f325;
                        p306 = p306 - tc;
                        p305 = p305 + tc;
                end
                327: begin
                        tc = f326;
                        p39 = p39 - tc;
                        p289 = p289 + tc;
                        p307 = p307 + tc;
                end
                328: begin
                        tc = f327;
                        p307 = p307 - tc;
                        p39 = p39 + tc;
                end
                329: begin
                        tc = f328;
                        p309 = p309 - tc;
                        p308 = p308 + tc;
                end
                330: begin
                        tc = f329;
                        p310 = p310 - tc;
                        p309 = p309 + tc;
                end
                331: begin
                        tc = f330;
                        p304 = p304 - tc;
                        p308 = p308 - tc;
                        p11 = p11 + tc;
                end
                332: begin
                        tc = f331;
                        p290 = p290 - tc;
                        p306 = p306 + tc;
                        p310 = p310 + tc;
                end
                333: begin
                        tc = f332;
                        p291 = p291 - tc;
                        p40 = p40 + tc;
                end
                334: begin
                        tc = f333;
                        p40 = p40 - tc;
                end
                335: begin
                        tc = f334;
                        p311 = p311 - tc;
                        p292 = p292 + tc;
                end
                336: begin
                        tc = f335;
                        p12 = p12 - tc;
                        p311 = p311 + tc;
                end
                337: begin
                        tc = f336;
                        p313 = p313 - tc;
                        p314 = p314 + tc;
                end
                338: begin
                        tc = f337;
                        p316 = p316 - tc;
                        p315 = p315 + tc;
                end
                339: begin
                        tc = f338;
                        p40 = p40 - tc;
                        p312 = p312 + tc;
                        p317 = p317 + tc;
                end
                340: begin
                        tc = f339;
                        p317 = p317 - tc;
                        p40 = p40 + tc;
                end
                341: begin
                        tc = f340;
                        p319 = p319 - tc;
                        p318 = p318 + tc;
                end
                342: begin
                        tc = f341;
                        p320 = p320 - tc;
                        p319 = p319 + tc;
                end
                343: begin
                        tc = f342;
                        p37 = p37 - tc;
                        p313 = p313 + tc;
                        p321 = p321 + tc;
                end
                344: begin
                        tc = f343;
                        p321 = p321 - tc;
                        p37 = p37 + tc;
                end
                345: begin
                        tc = f344;
                        p323 = p323 - tc;
                        p322 = p322 + tc;
                end
                346: begin
                        tc = f345;
                        p324 = p324 - tc;
                        p323 = p323 + tc;
                end
                347: begin
                        tc = f346;
                        p318 = p318 - tc;
                        p322 = p322 - tc;
                        p12 = p12 + tc;
                end
                348: begin
                        tc = f347;
                        p315 = p315 - tc;
                        p320 = p320 + tc;
                        p324 = p324 + tc;
                end
                349: begin
                        tc = f348;
                        p314 = p314 - tc;
                        p41 = p41 + tc;
                end
                350: begin
                        tc = f349;
                        p41 = p41 - tc;
                end
                351: begin
                        tc = f350;
                        p325 = p325 - tc;
                        p316 = p316 + tc;
                end
                352: begin
                        tc = f351;
                        p13 = p13 - tc;
                        p325 = p325 + tc;
                end
                353: begin
                        tc = f352;
                        p327 = p327 - tc;
                        p328 = p328 + tc;
                end
                354: begin
                        tc = f353;
                        p330 = p330 - tc;
                        p329 = p329 + tc;
                end
                355: begin
                        tc = f354;
                        p41 = p41 - tc;
                        p326 = p326 + tc;
                        p331 = p331 + tc;
                end
                356: begin
                        tc = f355;
                        p331 = p331 - tc;
                        p41 = p41 + tc;
                end
                357: begin
                        tc = f356;
                        p333 = p333 - tc;
                        p332 = p332 + tc;
                end
                358: begin
                        tc = f357;
                        p334 = p334 - tc;
                        p333 = p333 + tc;
                end
                359: begin
                        tc = f358;
                        p42 = p42 - tc;
                        p327 = p327 + tc;
                        p335 = p335 + tc;
                end
                360: begin
                        tc = f359;
                        p335 = p335 - tc;
                        p42 = p42 + tc;
                end
                361: begin
                        tc = f360;
                        p337 = p337 - tc;
                        p336 = p336 + tc;
                end
                362: begin
                        tc = f361;
                        p338 = p338 - tc;
                        p337 = p337 + tc;
                end
                363: begin
                        tc = f362;
                        p332 = p332 - tc;
                        p336 = p336 - tc;
                        p13 = p13 + tc;
                end
                364: begin
                        tc = f363;
                        p329 = p329 - tc;
                        p334 = p334 + tc;
                        p338 = p338 + tc;
                end
                365: begin
                        tc = f364;
                        p328 = p328 - tc;
                        p43 = p43 + tc;
                end
                366: begin
                        tc = f365;
                        p43 = p43 - tc;
                end
                367: begin
                        tc = f366;
                        p339 = p339 - tc;
                        p330 = p330 + tc;
                end
                368: begin
                        tc = f367;
                        p14 = p14 - tc;
                        p339 = p339 + tc;
                end
                default:;
        endcase
        led = ~p43[5:0];
end
end
endmodule