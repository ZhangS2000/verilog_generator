module sn(
	input clk,
	output reg [5:0] led
);
`define INH(place) ((place) == 0 ? 255 : 0)
reg [7:0] p0=0;
reg [7:0] p1=0;
reg [7:0] p2=0;
reg [7:0] p3=0;
reg [7:0] p4=0;
reg [7:0] p5=0;
reg [7:0] p6=0;
reg [7:0] p7=0;
reg [7:0] p8=0;
reg [7:0] p9=0;
reg [7:0] p10=0;
reg [7:0] p11=0;
reg [7:0] p12=0;
reg [7:0] p13=1;
reg [7:0] p14=2;
reg [7:0] p15=2;
reg [7:0] p16=2;
reg [7:0] p17=0;
reg [7:0] p18=0;
reg [7:0] p19=0;
reg [7:0] p20=0;
reg [7:0] p21=0;
reg [7:0] p22=0;
reg [7:0] p23=0;
reg [7:0] p24=0;
reg [7:0] p25=0;
reg [7:0] p26=0;
reg [7:0] p27=0;
reg [7:0] p28=0;
reg [7:0] p29=0;
reg [7:0] p30=0;
reg [7:0] p31=0;
reg [7:0] p32=0;
reg [7:0] p33=0;
reg [7:0] p34=0;
reg [7:0] p35=0;
reg [7:0] p36=0;
reg [7:0] p37=0;
reg [7:0] p38=0;
reg [7:0] p39=0;
reg [7:0] p40=0;
reg [7:0] p41=0;
reg [7:0] p42=0;
reg [7:0] p43=0;
reg [7:0] p44=0;
reg [7:0] p45=0;
reg [7:0] f[0:33];
reg [7:0] tf;
always @(posedge clk) begin
	f[0] = 255;
	f[0] = (f[0] > p0) ? p0 : f[0];
	f[0] = (f[0] > p15) ? p15 : f[0];
	f[1] = 255;
	f[1] = (f[1] > p2) ? p2 : f[1];
	f[1] = (f[1] > p10) ? p10 : f[1];
	f[1] = (f[1] > p11) ? p11 : f[1];
	f[2] = 255;
	f[2] = (f[2] > p3) ? p3 : f[2];
	f[2] = (f[2] > p7) ? p7 : f[2];
	f[2] = (f[2] > p11) ? p11 : f[2];
	f[3] = 255;
	f[3] = (f[3] > p2) ? p2 : f[3];
	f[3] = (f[3] > p8) ? p8 : f[3];
	f[3] = (f[3] > p10) ? p10 : f[3];
	f[4] = 255;
	f[4] = (f[4] > p4) ? p4 : f[4];
	f[5] = 255;
	f[5] = (f[5] > p6) ? p6 : f[5];
	f[6] = 255;
	f[6] = (f[6] > p3) ? p3 : f[6];
	f[6] = (f[6] > p7) ? p7 : f[6];
	f[6] = (f[6] > p8) ? p8 : f[6];
	f[7] = 255;
	f[7] = (f[7] > p4) ? p4 : f[7];
	f[7] = (f[7] > p10) ? p10 : f[7];
	f[7] = (f[7] > p15) ? p15 : f[7];
	f[8] = 255;
	f[8] = (f[8] > p6) ? p6 : f[8];
	f[8] = (f[8] > p7) ? p7 : f[8];
	f[8] = (f[8] > p9) ? p9 : f[8];
	f[8] = (f[8] > p16) ? p16 : f[8];
	f[9] = 255;
	f[9] = (f[9] > p1) ? p1 : f[9];
	f[9] = (f[9] > p6) ? p6 : f[9];
	f[9] = (f[9] > p10) ? p10 : f[9];
	f[9] = (f[9] > p16) ? p16 : f[9];
	f[10] = 255;
	f[10] = (f[10] > p4) ? p4 : f[10];
	f[10] = (f[10] > p7) ? p7 : f[10];
	f[10] = (f[10] > p14) ? p14 : f[10];
	f[11] = 255;
	f[11] = (f[11] > p13) ? p13 : f[11];
	f[11] = (f[11] > p14) ? p14 : f[11];
	f[12] = 255;
	f[12] = (f[12] > p12) ? p12 : f[12];
	f[12] = (f[12] > p19) ? p19 : f[12];
	f[13] = 255;
	f[13] = (f[13] > p5) ? p5 : f[13];
	f[13] = (f[13] > p17) ? p17 : f[13];
	f[14] = 255;
	f[14] = (f[14] > p5) ? p5 : f[14];
	f[14] = (f[14] > p18) ? p18 : f[14];
	f[15] = 255;
	f[15] = (f[15] > p20) ? p20 : f[15];
	f[15] = (f[15] > p35) ? p35 : f[15];
	f[16] = 255;
	f[16] = (f[16] > p22) ? p22 : f[16];
	f[16] = (f[16] > p30) ? p30 : f[16];
	f[16] = (f[16] > p31) ? p31 : f[16];
	f[17] = 255;
	f[17] = (f[17] > p23) ? p23 : f[17];
	f[17] = (f[17] > p27) ? p27 : f[17];
	f[17] = (f[17] > p31) ? p31 : f[17];
	f[18] = 255;
	f[18] = (f[18] > p22) ? p22 : f[18];
	f[18] = (f[18] > p28) ? p28 : f[18];
	f[18] = (f[18] > p30) ? p30 : f[18];
	f[19] = 255;
	f[19] = (f[19] > p24) ? p24 : f[19];
	f[20] = 255;
	f[20] = (f[20] > p26) ? p26 : f[20];
	f[21] = 255;
	f[21] = (f[21] > p23) ? p23 : f[21];
	f[21] = (f[21] > p27) ? p27 : f[21];
	f[21] = (f[21] > p28) ? p28 : f[21];
	f[22] = 255;
	f[22] = (f[22] > p24) ? p24 : f[22];
	f[22] = (f[22] > p30) ? p30 : f[22];
	f[22] = (f[22] > p35) ? p35 : f[22];
	f[23] = 255;
	f[23] = (f[23] > p26) ? p26 : f[23];
	f[23] = (f[23] > p27) ? p27 : f[23];
	f[23] = (f[23] > p29) ? p29 : f[23];
	f[23] = (f[23] > p36) ? p36 : f[23];
	f[24] = 255;
	f[24] = (f[24] > p21) ? p21 : f[24];
	f[24] = (f[24] > p26) ? p26 : f[24];
	f[24] = (f[24] > p30) ? p30 : f[24];
	f[24] = (f[24] > p36) ? p36 : f[24];
	f[25] = 255;
	f[25] = (f[25] > p24) ? p24 : f[25];
	f[25] = (f[25] > p27) ? p27 : f[25];
	f[25] = (f[25] > p34) ? p34 : f[25];
	f[26] = 255;
	f[26] = (f[26] > p33) ? p33 : f[26];
	f[26] = (f[26] > p34) ? p34 : f[26];
	f[27] = 255;
	f[27] = (f[27] > p32) ? p32 : f[27];
	f[27] = (f[27] > p41) ? p41 : f[27];
	f[28] = 255;
	f[28] = (f[28] > p14) ? p14 : f[28];
	f[28] = (f[28] > p37) ? p37 : f[28];
	f[29] = 255;
	f[29] = (f[29] > p15) ? p15 : f[29];
	f[29] = (f[29] > p25) ? p25 : f[29];
	f[29] = (f[29] > p38) ? p38 : f[29];
	f[30] = 255;
	f[30] = (f[30] > p8) ? p8 : f[30];
	f[30] = (f[30] > p10) ? p10 : f[30];
	f[30] = (f[30] > p39) ? p39 : f[30];
	f[31] = 255;
	f[31] = (f[31] > p10) ? p10 : f[31];
	f[31] = (f[31] > p11) ? p11 : f[31];
	f[31] = (f[31] > p39) ? p39 : f[31];
	f[32] = 255;
	f[32] = (f[32] > p7) ? p7 : f[32];
	f[32] = (f[32] > p8) ? p8 : f[32];
	f[32] = (f[32] > p40) ? p40 : f[32];
	f[33] = 255;
	f[33] = (f[33] > p7) ? p7 : f[33];
	f[33] = (f[33] > p11) ? p11 : f[33];
	f[33] = (f[33] > p40) ? p40 : f[33];
    if(f[0]>0) tf = 0;
    else if(f[1]>0) tf = 1;
    else if(f[2]>0) tf = 2;
    else if(f[3]>0) tf = 3;
    else if(f[6]>0) tf = 6;
    else if(f[7]>0) tf = 7;
    else if(f[8]>0) tf = 8;
    else if(f[9]>0) tf = 9;
    else if(f[10]>0) tf = 10;
    else if(f[11]>0) tf = 11;
    else if(f[12]>0) tf = 12;
    else if(f[13]>0) tf = 13;
    else if(f[14]>0) tf = 14;
    else if(f[15]>0) tf = 15;
    else if(f[16]>0) tf = 16;
    else if(f[17]>0) tf = 17;
    else if(f[18]>0) tf = 18;
    else if(f[21]>0) tf = 21;
    else if(f[22]>0) tf = 22;
    else if(f[23]>0) tf = 23;
    else if(f[24]>0) tf = 24;
    else if(f[25]>0) tf = 25;
    else if(f[26]>0) tf = 26;
    else if(f[27]>0) tf = 27;
    else if(f[28]>0) tf = 28;
    else if(f[29]>0) tf = 29;
    else if(f[30]>0) tf = 30;
    else if(f[31]>0) tf = 31;
    else if(f[32]>0) tf = 32;
    else if(f[33]>0) tf = 33;
    else if(f[4]>0) tf = 4;
    else if(f[5]>0) tf = 5;
    else if(f[19]>0) tf = 19;
    else if(f[20]>0) tf = 20;
    else tf = 34;
	case(tf)
		0: begin
			p0 = p0 - f[0];
			p15 = p15 - f[0];
			p1 = p1 + f[0];
			p2 = p2 + f[0];
			p4 = p4 + f[0];
			p10 = p10 + f[0];
			p34 = p34 + f[0];
			p35 = p35 + f[0];
			p36 = p36 + f[0];
		end
		1: begin
			p2 = p2 - f[1];
			p10 = p10 - f[1];
			p11 = p11 - f[1];
			p3 = p3 + f[1];
			p4 = p4 + f[1];
			p7 = p7 + f[1];
		end
		2: begin
			p3 = p3 - f[2];
			p7 = p7 - f[2];
			p11 = p11 - f[2];
			p33 = p33 + f[2];
		end
		3: begin
			p2 = p2 - f[3];
			p8 = p8 - f[3];
			p10 = p10 - f[3];
			p0 = p0 + f[3];
		end
		4: begin
			p4 = p4 - f[6];
			p6 = p6 + f[6];
		end
		5: begin
			p6 = p6 - f[7];
			p12 = p12 + f[7];
			p17 = p17 + f[7];
		end
		6: begin
			p3 = p3 - f[8];
			p7 = p7 - f[8];
			p8 = p8 - f[8];
			p13 = p13 + f[8];
		end
		7: begin
			p4 = p4 - f[9];
			p10 = p10 - f[9];
			p15 = p15 - f[9];
			p8 = p8 + f[9];
			p10 = p10 + f[9];
			p15 = p15 + f[9];
		end
		8: begin
			p6 = p6 - f[10];
			p7 = p7 - f[10];
			p9 = p9 - f[10];
			p16 = p16 - f[10];
			p5 = p5 + f[10];
			p6 = p6 + f[10];
			p7 = p7 + f[10];
			p14 = p14 + f[10];
		end
		9: begin
			p1 = p1 - f[11];
			p6 = p6 - f[11];
			p10 = p10 - f[11];
			p16 = p16 - f[11];
			p5 = p5 + f[11];
			p6 = p6 + f[11];
			p10 = p10 + f[11];
			p15 = p15 + f[11];
		end
		10: begin
			p4 = p4 - f[12];
			p7 = p7 - f[12];
			p14 = p14 - f[12];
			p7 = p7 + f[12];
			p8 = p8 + f[12];
			p14 = p14 + f[12];
		end
		11: begin
			p13 = p13 - f[13];
			p14 = p14 - f[13];
			p0 = p0 + f[13];
			p9 = p9 + f[13];
		end
		12: begin
			p12 = p12 - f[14];
			p19 = p19 - f[14];
			p11 = p11 + f[14];
		end
		13: begin
			p5 = p5 - f[15];
			p17 = p17 - f[15];
			p16 = p16 + f[15];
			p18 = p18 + f[15];
		end
		14: begin
			p5 = p5 - f[16];
			p18 = p18 - f[16];
			p16 = p16 + f[16];
			p19 = p19 + f[16];
		end
		15: begin
			p20 = p20 - f[17];
			p35 = p35 - f[17];
			p21 = p21 + f[17];
			p22 = p22 + f[17];
			p24 = p24 + f[17];
			p30 = p30 + f[17];
			p43 = p43 + f[17];
			p44 = p44 + f[17];
			p45 = p45 + f[17];
		end
		16: begin
			p22 = p22 - f[18];
			p30 = p30 - f[18];
			p31 = p31 - f[18];
			p23 = p23 + f[18];
			p24 = p24 + f[18];
			p27 = p27 + f[18];
		end
		17: begin
			p23 = p23 - f[21];
			p27 = p27 - f[21];
			p31 = p31 - f[21];
			p42 = p42 + f[21];
		end
		18: begin
			p22 = p22 - f[22];
			p28 = p28 - f[22];
			p30 = p30 - f[22];
			p20 = p20 + f[22];
		end
		19: begin
			p24 = p24 - f[23];
			p26 = p26 + f[23];
		end
		20: begin
			p26 = p26 - f[24];
			p32 = p32 + f[24];
			p37 = p37 + f[24];
		end
		21: begin
			p23 = p23 - f[25];
			p27 = p27 - f[25];
			p28 = p28 - f[25];
			p33 = p33 + f[25];
		end
		22: begin
			p24 = p24 - f[26];
			p30 = p30 - f[26];
			p35 = p35 - f[26];
			p28 = p28 + f[26];
			p30 = p30 + f[26];
			p35 = p35 + f[26];
		end
		23: begin
			p26 = p26 - f[27];
			p27 = p27 - f[27];
			p29 = p29 - f[27];
			p36 = p36 - f[27];
			p25 = p25 + f[27];
			p26 = p26 + f[27];
			p27 = p27 + f[27];
			p34 = p34 + f[27];
		end
		24: begin
			p21 = p21 - f[28];
			p26 = p26 - f[28];
			p30 = p30 - f[28];
			p36 = p36 - f[28];
			p25 = p25 + f[28];
			p26 = p26 + f[28];
			p30 = p30 + f[28];
			p35 = p35 + f[28];
		end
		25: begin
			p24 = p24 - f[29];
			p27 = p27 - f[29];
			p34 = p34 - f[29];
			p27 = p27 + f[29];
			p28 = p28 + f[29];
			p34 = p34 + f[29];
		end
		26: begin
			p33 = p33 - f[30];
			p34 = p34 - f[30];
			p20 = p20 + f[30];
			p29 = p29 + f[30];
		end
		27: begin
			p32 = p32 - f[31];
			p41 = p41 - f[31];
			p31 = p31 + f[31];
		end
		28: begin
			p14 = p14 - f[32];
			p37 = p37 - f[32];
			p9 = p9 + f[32];
			p38 = p38 + f[32];
		end
		29: begin
			p15 = p15 - f[33];
			p25 = p25 - f[33];
			p38 = p38 - f[33];
			p1 = p1 + f[33];
			p4 = p4 + f[33];
			p10 = p10 + f[33];
			p36 = p36 + f[33];
			p39 = p39 + f[33];
		end
		30: begin
			p8 = p8 - f[4];
			p10 = p10 - f[4];
			p39 = p39 - f[4];
			p38 = p38 + f[4];
		end
		31: begin
			p10 = p10 - f[5];
			p11 = p11 - f[5];
			p39 = p39 - f[5];
			p4 = p4 + f[5];
			p7 = p7 + f[5];
			p40 = p40 + f[5];
		end
		32: begin
			p7 = p7 - f[19];
			p8 = p8 - f[19];
			p40 = p40 - f[19];
			p37 = p37 + f[19];
		end
		33: begin
			p7 = p7 - f[20];
			p11 = p11 - f[20];
			p40 = p40 - f[20];
			p41 = p41 + f[20];
		end
		default:;
	endcase
	led = ~p45[5:0];
end
endmodule