module sn(
        input clk,
        output reg [5:0] led
);

`define C0 8'b00000000
`define C1 8'b00000001
`define C2 8'b00000010
`define C5 8'b00000101
`define C8 8'b00001000
`define C255 8'b11111111

`define INH( x ) (((x) == `C0) ? `C255 : `C0)

reg [7:0] p [116:0]= {`C0,`C1,`C1,`C1,`C1,`C1,`C8,`C2,`C0,`C2,`C0,`C5,`C2,`C0,`C0,`C1,`C0,`C0,`C0,`C1,`C0,`C1,`C1,`C1,`C0,`C1,`C0,`C1,`C1,`C0,`C1,`C1,`C0,`C1,`C1,`C1,`C0,`C1,`C1,`C1,`C1,`C0,`C0,`C1,`C0,`C1,`C1,`C1,`C0,`C1,`C0,`C1,`C1,`C0,`C1,`C1,`C0,`C1,`C1,`C1,`C0,`C1,`C1,`C1,`C1,`C0,`C0,`C1,`C0,`C1,`C1,`C1,`C0,`C1,`C0,`C1,`C1,`C0,`C1,`C1,`C0,`C1,`C1,`C1,`C0,`C1,`C1,`C1,`C1,`C0,`C0,`C0,`C1,`C1,`C0,`C1,`C1,`C1,`C0,`C1,`C1,`C1,`C1,`C0,`C0,`C0,`C1,`C1,`C0,`C1,`C1,`C1,`C0,`C1,`C1,`C1,`C1};
reg [7:0] y [0: 123];
//initial
//begin
//p[0]=`C0; p[1]=`C1; p[2]=`C1; p[3]=`C1; p[4]=`C1; p[5]=`C1; p[6]=`C8; p[7]=`C2; p[8]=`C0; p[9]=`C2; 
//p[10]=`C0; p[11]=`C5; p[12]=`C2; p[13]=`C0; p[14]=`C0; p[15]=`C1; p[16]=`C0; p[17]=`C0; p[18]=`C0; p[19]=`C1; 
//p[20]=`C0; p[21]=`C1; p[22]=`C1; p[23]=`C1; p[24]=`C0; p[25]=`C1; p[26]=`C0; p[27]=`C1; p[28]=`C1; p[29]=`C0; 
//p[30]=`C1; p[31]=`C1; p[32]=`C0; p[33]=`C1; p[34]=`C1; p[35]=`C1; p[36]=`C0; p[37]=`C1; p[38]=`C1; p[39]=`C1; 
//p[40]=`C1; p[41]=`C0; p[42]=`C0; p[43]=`C1; p[44]=`C0; p[45]=`C1; p[46]=`C1; p[47]=`C1; p[48]=`C0; p[49]=`C1; 
//p[50]=`C0; p[51]=`C1; p[52]=`C1; p[53]=`C0; p[54]=`C1; p[55]=`C1; p[56]=`C0; p[57]=`C1; p[58]=`C1; p[59]=`C1; 
//p[60]=`C0; p[61]=`C1; p[62]=`C1; p[63]=`C1; p[64]=`C1; p[65]=`C0; p[66]=`C0; p[67]=`C1; p[68]=`C0; p[69]=`C1; 
//p[70]=`C1; p[71]=`C1; p[72]=`C0; p[73]=`C1; p[74]=`C0; p[75]=`C1; p[76]=`C1; p[77]=`C0; p[78]=`C1; p[79]=`C1; 
//p[80]=`C0; p[81]=`C1; p[82]=`C1; p[83]=`C1; p[84]=`C0; p[85]=`C1; p[86]=`C1; p[87]=`C1; p[88]=`C1; p[89]=`C0; 
//p[90]=`C0; p[91]=`C0; p[92]=`C1; p[93]=`C1; p[94]=`C0; p[95]=`C1; p[96]=`C1; p[97]=`C1; p[98]=`C0; p[99]=`C1; 
//p[100]=`C1; p[101]=`C1; p[102]=`C1; p[103]=`C0; p[104]=`C0; p[105]=`C0; p[106]=`C1; p[107]=`C1; p[108]=`C0; p[109]=`C1; 
//p[110]=`C1; p[111]=`C1; p[112]=`C0; p[113]=`C1; p[114]=`C1; p[115]=`C1; p[116]=`C1; 
//end


always @(posedge clk) begin
        y[0] = `C255;
        y[0] = (y[0] > `INH(p[19])) ? `INH(p[19]) : y[0];
        y[0] = (y[0] > p[22]) ? p[22] : y[0];
        y[1] = `C255;
        y[1] = (y[1] > `INH(p[43])) ? `INH(p[43]) : y[1];
        y[1] = (y[1] > p[46]) ? p[46] : y[1];
        y[2] = `C255;
        y[2] = (y[2] > `INH(p[67])) ? `INH(p[67]) : y[2];
        y[2] = (y[2] > p[70]) ? p[70] : y[2];
        y[3] = `C255;
        y[3] = (y[3] > p[89]) ? p[89] : y[3];
        y[3] = (y[3] > `INH(p[92])) ? `INH(p[92]) : y[3];
        y[4] = `C255;
        y[4] = (y[4] > p[103]) ? p[103] : y[4];
        y[4] = (y[4] > `INH(p[106])) ? `INH(p[106]) : y[4];
        y[5] = `C255;
        y[5] = (y[5] > `INH(p[18])) ? `INH(p[18]) : y[5];
        y[5] = (y[5] > `INH(p[19])) ? `INH(p[19]) : y[5];
        y[5] = (y[5] > p[23]) ? p[23] : y[5];
        y[6] = `C255;
        y[6] = (y[6] > p[17]) ? p[17] : y[6];
        y[6] = (y[6] > `INH(p[23])) ? `INH(p[23]) : y[6];
        y[7] = `C255;
        y[7] = (y[7] > p[21]) ? p[21] : y[7];
        y[7] = (y[7] > `INH(p[23])) ? `INH(p[23]) : y[7];
        y[8] = `C255;
        y[8] = (y[8] > p[18/2]) ? p[18/2] : y[8];
        y[8] = (y[8] > `INH(p[22])) ? `INH(p[22]) : y[8];
        y[9] = `C255;
        y[9] = (y[9] > `INH(p[22])) ? `INH(p[22]) : y[9];
        y[9] = (y[9] > p[25]) ? p[25] : y[9];
        y[10] = `C255;
        y[10] = (y[10] > p[18]) ? p[18] : y[10];
        y[10] = (y[10] > `INH(p[25])) ? `INH(p[25]) : y[10];
        y[10] = (y[10] > p[27]) ? p[27] : y[10];
        y[11] = `C255;
        y[11] = (y[11] > `INH(p[25])) ? `INH(p[25]) : y[11];
        y[11] = (y[11] > p[28]) ? p[28] : y[11];
        y[12] = `C255;
        y[12] = (y[12] > p[17]) ? p[17] : y[12];
        y[12] = (y[12] > `INH(p[27])) ? `INH(p[27]) : y[12];
        y[12] = (y[12] > `INH(p[28])) ? `INH(p[28]) : y[12];
        y[13] = `C255;
        y[13] = (y[13] > p[17]) ? p[17] : y[13];
        y[13] = (y[13] > `INH(p[26])) ? `INH(p[26]) : y[13];
        y[13] = (y[13] > `INH(p[28])) ? `INH(p[28]) : y[13];
        y[14] = `C255;
        y[14] = (y[14] > `INH(p[28])) ? `INH(p[28]) : y[14];
        y[14] = (y[14] > p[30]) ? p[30] : y[14];
        y[15] = `C255;
        y[15] = (y[15] > p[24]) ? p[24] : y[15];
        y[15] = (y[15] > `INH(p[30])) ? `INH(p[30]) : y[15];
        y[16] = `C255;
        y[16] = (y[16] > `INH(p[30])) ? `INH(p[30]) : y[16];
        y[16] = (y[16] > p[31]) ? p[31] : y[16];
        y[17] = `C255;
        y[17] = (y[17] > p[29]) ? p[29] : y[17];
        y[17] = (y[17] > `INH(p[31])) ? `INH(p[31]) : y[17];
        y[18] = `C255;
        y[18] = (y[18] > p[19]) ? p[19] : y[18];
        y[18] = (y[18] > p[26]) ? p[26] : y[18];
        y[18] = (y[18] > `INH(p[27])) ? `INH(p[27]) : y[18];
        y[18] = (y[18] > `INH(p[31])) ? `INH(p[31]) : y[18];
        y[19] = `C255;
        y[19] = (y[19] > p[19]) ? p[19] : y[19];
        y[19] = (y[19] > `INH(p[26])) ? `INH(p[26]) : y[19];
        y[19] = (y[19] > `INH(p[31])) ? `INH(p[31]) : y[19];
        y[20] = `C255;
        y[20] = (y[20] > p[6]) ? p[6] : y[20];
        y[20] = (y[20] > `INH(p[33])) ? `INH(p[33]) : y[20];
        y[21] = `C255;
        y[21] = (y[21] > p[32]) ? p[32] : y[21];
        y[21] = (y[21] > `INH(p[34])) ? `INH(p[34]) : y[21];
        y[22] = `C255;
        y[22] = (y[22] > `INH(p[6])) ? `INH(p[6]) : y[22];
        y[22] = (y[22] > `INH(p[33])) ? `INH(p[33]) : y[22];
        y[22] = (y[22] > p[34]) ? p[34] : y[22];
        y[23] = `C255;
        y[23] = (y[23] > `INH(p[32])) ? `INH(p[32]) : y[23];
        y[23] = (y[23] > `INH(p[34])) ? `INH(p[34]) : y[23];
        y[23] = (y[23] > p[35]) ? p[35] : y[23];
        y[24] = `C255;
        y[24] = (y[24] > p[7]) ? p[7] : y[24];
        y[24] = (y[24] > `INH(p[37])) ? `INH(p[37]) : y[24];
        y[25] = `C255;
        y[25] = (y[25] > p[36]) ? p[36] : y[25];
        y[25] = (y[25] > `INH(p[38])) ? `INH(p[38]) : y[25];
        y[26] = `C255;
        y[26] = (y[26] > `INH(p[7])) ? `INH(p[7]) : y[26];
        y[26] = (y[26] > `INH(p[37])) ? `INH(p[37]) : y[26];
        y[26] = (y[26] > p[38]) ? p[38] : y[26];
        y[27] = `C255;
        y[27] = (y[27] > `INH(p[36])) ? `INH(p[36]) : y[27];
        y[27] = (y[27] > `INH(p[38])) ? `INH(p[38]) : y[27];
        y[27] = (y[27] > p[39]) ? p[39] : y[27];
        y[28] = `C255;
        y[28] = (y[28] > `INH(p[0])) ? `INH(p[0]) : y[28];
        y[28] = (y[28] > p[33]) ? p[33] : y[28];
        y[28] = (y[28] > p[37]) ? p[37] : y[28];
        y[29] = `C255;
        y[29] = (y[29] > p[19]) ? p[19] : y[29];
        y[29] = (y[29] > `INH(p[35])) ? `INH(p[35]) : y[29];
        y[29] = (y[29] > `INH(p[39])) ? `INH(p[39]) : y[29];
        y[30] = `C255;
        y[30] = (y[30] > p[20]) ? p[20] : y[30];
        y[30] = (y[30] > `INH(p[40])) ? `INH(p[40]) : y[30];
        y[31] = `C255;
        y[31] = (y[31] > p[8]) ? p[8] : y[31];
        y[31] = (y[31] > `INH(p[21])) ? `INH(p[21]) : y[31];
        y[32] = `C255;
        y[32] = (y[32] > `INH(p[8])) ? `INH(p[8]) : y[32];
        y[32] = (y[32] > `INH(p[21])) ? `INH(p[21]) : y[32];
        y[32] = (y[32] > p[40]) ? p[40] : y[32];
        y[33] = `C255;
        y[33] = (y[33] > p[1]) ? p[1] : y[33];
        y[33] = (y[33] > `INH(p[20])) ? `INH(p[20]) : y[33];
        y[33] = (y[33] > `INH(p[40])) ? `INH(p[40]) : y[33];
        y[34] = `C255;
        y[34] = (y[34] > `INH(p[42])) ? `INH(p[42]) : y[34];
        y[34] = (y[34] > `INH(p[43])) ? `INH(p[43]) : y[34];
        y[34] = (y[34] > p[47]) ? p[47] : y[34];
        y[35] = `C255;
        y[35] = (y[35] > p[41]) ? p[41] : y[35];
        y[35] = (y[35] > `INH(p[47])) ? `INH(p[47]) : y[35];
        y[36] = `C255;
        y[36] = (y[36] > p[45]) ? p[45] : y[36];
        y[36] = (y[36] > `INH(p[47])) ? `INH(p[47]) : y[36];
        y[37] = `C255;
        y[37] = (y[37] > p[42/2]) ? p[42/2] : y[37];
        y[37] = (y[37] > `INH(p[46])) ? `INH(p[46]) : y[37];
        y[38] = `C255;
        y[38] = (y[38] > `INH(p[46])) ? `INH(p[46]) : y[38];
        y[38] = (y[38] > p[49]) ? p[49] : y[38];
        y[39] = `C255;
        y[39] = (y[39] > p[42]) ? p[42] : y[39];
        y[39] = (y[39] > `INH(p[49])) ? `INH(p[49]) : y[39];
        y[39] = (y[39] > p[51]) ? p[51] : y[39];
        y[40] = `C255;
        y[40] = (y[40] > `INH(p[49])) ? `INH(p[49]) : y[40];
        y[40] = (y[40] > p[52]) ? p[52] : y[40];
        y[41] = `C255;
        y[41] = (y[41] > p[41]) ? p[41] : y[41];
        y[41] = (y[41] > `INH(p[51])) ? `INH(p[51]) : y[41];
        y[41] = (y[41] > `INH(p[52])) ? `INH(p[52]) : y[41];
        y[42] = `C255;
        y[42] = (y[42] > p[41]) ? p[41] : y[42];
        y[42] = (y[42] > `INH(p[50])) ? `INH(p[50]) : y[42];
        y[42] = (y[42] > `INH(p[52])) ? `INH(p[52]) : y[42];
        y[43] = `C255;
        y[43] = (y[43] > `INH(p[52])) ? `INH(p[52]) : y[43];
        y[43] = (y[43] > p[54]) ? p[54] : y[43];
        y[44] = `C255;
        y[44] = (y[44] > p[48]) ? p[48] : y[44];
        y[44] = (y[44] > `INH(p[54])) ? `INH(p[54]) : y[44];
        y[45] = `C255;
        y[45] = (y[45] > `INH(p[54])) ? `INH(p[54]) : y[45];
        y[45] = (y[45] > p[55]) ? p[55] : y[45];
        y[46] = `C255;
        y[46] = (y[46] > p[53]) ? p[53] : y[46];
        y[46] = (y[46] > `INH(p[55])) ? `INH(p[55]) : y[46];
        y[47] = `C255;
        y[47] = (y[47] > p[43]) ? p[43] : y[47];
        y[47] = (y[47] > p[50]) ? p[50] : y[47];
        y[47] = (y[47] > `INH(p[51])) ? `INH(p[51]) : y[47];
        y[47] = (y[47] > `INH(p[55])) ? `INH(p[55]) : y[47];
        y[48] = `C255;
        y[48] = (y[48] > p[43]) ? p[43] : y[48];
        y[48] = (y[48] > `INH(p[50])) ? `INH(p[50]) : y[48];
        y[48] = (y[48] > `INH(p[55])) ? `INH(p[55]) : y[48];
        y[49] = `C255;
        y[49] = (y[49] > p[8]) ? p[8] : y[49];
        y[49] = (y[49] > `INH(p[57])) ? `INH(p[57]) : y[49];
        y[50] = `C255;
        y[50] = (y[50] > p[56]) ? p[56] : y[50];
        y[50] = (y[50] > `INH(p[58])) ? `INH(p[58]) : y[50];
        y[51] = `C255;
        y[51] = (y[51] > `INH(p[8])) ? `INH(p[8]) : y[51];
        y[51] = (y[51] > `INH(p[57])) ? `INH(p[57]) : y[51];
        y[51] = (y[51] > p[58]) ? p[58] : y[51];
        y[52] = `C255;
        y[52] = (y[52] > `INH(p[56])) ? `INH(p[56]) : y[52];
        y[52] = (y[52] > `INH(p[58])) ? `INH(p[58]) : y[52];
        y[52] = (y[52] > p[59]) ? p[59] : y[52];
        y[53] = `C255;
        y[53] = (y[53] > p[9]) ? p[9] : y[53];
        y[53] = (y[53] > `INH(p[61])) ? `INH(p[61]) : y[53];
        y[54] = `C255;
        y[54] = (y[54] > p[60]) ? p[60] : y[54];
        y[54] = (y[54] > `INH(p[62])) ? `INH(p[62]) : y[54];
        y[55] = `C255;
        y[55] = (y[55] > `INH(p[9])) ? `INH(p[9]) : y[55];
        y[55] = (y[55] > `INH(p[61])) ? `INH(p[61]) : y[55];
        y[55] = (y[55] > p[62]) ? p[62] : y[55];
        y[56] = `C255;
        y[56] = (y[56] > `INH(p[60])) ? `INH(p[60]) : y[56];
        y[56] = (y[56] > `INH(p[62])) ? `INH(p[62]) : y[56];
        y[56] = (y[56] > p[63]) ? p[63] : y[56];
        y[57] = `C255;
        y[57] = (y[57] > `INH(p[1])) ? `INH(p[1]) : y[57];
        y[57] = (y[57] > p[57]) ? p[57] : y[57];
        y[57] = (y[57] > p[61]) ? p[61] : y[57];
        y[58] = `C255;
        y[58] = (y[58] > p[43]) ? p[43] : y[58];
        y[58] = (y[58] > `INH(p[59])) ? `INH(p[59]) : y[58];
        y[58] = (y[58] > `INH(p[63])) ? `INH(p[63]) : y[58];
        y[59] = `C255;
        y[59] = (y[59] > p[44]) ? p[44] : y[59];
        y[59] = (y[59] > `INH(p[64])) ? `INH(p[64]) : y[59];
        y[60] = `C255;
        y[60] = (y[60] > p[10]) ? p[10] : y[60];
        y[60] = (y[60] > `INH(p[45])) ? `INH(p[45]) : y[60];
        y[61] = `C255;
        y[61] = (y[61] > `INH(p[10])) ? `INH(p[10]) : y[61];
        y[61] = (y[61] > `INH(p[45])) ? `INH(p[45]) : y[61];
        y[61] = (y[61] > p[64]) ? p[64] : y[61];
        y[62] = `C255;
        y[62] = (y[62] > p[2]) ? p[2] : y[62];
        y[62] = (y[62] > `INH(p[44])) ? `INH(p[44]) : y[62];
        y[62] = (y[62] > `INH(p[64])) ? `INH(p[64]) : y[62];
        y[63] = `C255;
        y[63] = (y[63] > `INH(p[66])) ? `INH(p[66]) : y[63];
        y[63] = (y[63] > `INH(p[67])) ? `INH(p[67]) : y[63];
        y[63] = (y[63] > p[71]) ? p[71] : y[63];
        y[64] = `C255;
        y[64] = (y[64] > p[65]) ? p[65] : y[64];
        y[64] = (y[64] > `INH(p[71])) ? `INH(p[71]) : y[64];
        y[65] = `C255;
        y[65] = (y[65] > p[69]) ? p[69] : y[65];
        y[65] = (y[65] > `INH(p[71])) ? `INH(p[71]) : y[65];
        y[66] = `C255;
        y[66] = (y[66] > p[66/2]) ? p[66/2] : y[66];
        y[66] = (y[66] > `INH(p[70])) ? `INH(p[70]) : y[66];
        y[67] = `C255;
        y[67] = (y[67] > `INH(p[70])) ? `INH(p[70]) : y[67];
        y[67] = (y[67] > p[73]) ? p[73] : y[67];
        y[68] = `C255;
        y[68] = (y[68] > p[66]) ? p[66] : y[68];
        y[68] = (y[68] > `INH(p[73])) ? `INH(p[73]) : y[68];
        y[68] = (y[68] > p[75]) ? p[75] : y[68];
        y[69] = `C255;
        y[69] = (y[69] > `INH(p[73])) ? `INH(p[73]) : y[69];
        y[69] = (y[69] > p[76]) ? p[76] : y[69];
        y[70] = `C255;
        y[70] = (y[70] > p[65]) ? p[65] : y[70];
        y[70] = (y[70] > `INH(p[75])) ? `INH(p[75]) : y[70];
        y[70] = (y[70] > `INH(p[76])) ? `INH(p[76]) : y[70];
        y[71] = `C255;
        y[71] = (y[71] > p[65]) ? p[65] : y[71];
        y[71] = (y[71] > `INH(p[74])) ? `INH(p[74]) : y[71];
        y[71] = (y[71] > `INH(p[76])) ? `INH(p[76]) : y[71];
        y[72] = `C255;
        y[72] = (y[72] > `INH(p[76])) ? `INH(p[76]) : y[72];
        y[72] = (y[72] > p[78]) ? p[78] : y[72];
        y[73] = `C255;
        y[73] = (y[73] > p[72]) ? p[72] : y[73];
        y[73] = (y[73] > `INH(p[78])) ? `INH(p[78]) : y[73];
        y[74] = `C255;
        y[74] = (y[74] > `INH(p[78])) ? `INH(p[78]) : y[74];
        y[74] = (y[74] > p[79]) ? p[79] : y[74];
        y[75] = `C255;
        y[75] = (y[75] > p[77]) ? p[77] : y[75];
        y[75] = (y[75] > `INH(p[79])) ? `INH(p[79]) : y[75];
        y[76] = `C255;
        y[76] = (y[76] > p[67]) ? p[67] : y[76];
        y[76] = (y[76] > p[74]) ? p[74] : y[76];
        y[76] = (y[76] > `INH(p[75])) ? `INH(p[75]) : y[76];
        y[76] = (y[76] > `INH(p[79])) ? `INH(p[79]) : y[76];
        y[77] = `C255;
        y[77] = (y[77] > p[67]) ? p[67] : y[77];
        y[77] = (y[77] > `INH(p[74])) ? `INH(p[74]) : y[77];
        y[77] = (y[77] > `INH(p[79])) ? `INH(p[79]) : y[77];
        y[78] = `C255;
        y[78] = (y[78] > p[11]) ? p[11] : y[78];
        y[78] = (y[78] > `INH(p[81])) ? `INH(p[81]) : y[78];
        y[79] = `C255;
        y[79] = (y[79] > p[80]) ? p[80] : y[79];
        y[79] = (y[79] > `INH(p[82])) ? `INH(p[82]) : y[79];
        y[80] = `C255;
        y[80] = (y[80] > `INH(p[11])) ? `INH(p[11]) : y[80];
        y[80] = (y[80] > `INH(p[81])) ? `INH(p[81]) : y[80];
        y[80] = (y[80] > p[82]) ? p[82] : y[80];
        y[81] = `C255;
        y[81] = (y[81] > `INH(p[80])) ? `INH(p[80]) : y[81];
        y[81] = (y[81] > `INH(p[82])) ? `INH(p[82]) : y[81];
        y[81] = (y[81] > p[83]) ? p[83] : y[81];
        y[82] = `C255;
        y[82] = (y[82] > p[12]) ? p[12] : y[82];
        y[82] = (y[82] > `INH(p[85])) ? `INH(p[85]) : y[82];
        y[83] = `C255;
        y[83] = (y[83] > p[84]) ? p[84] : y[83];
        y[83] = (y[83] > `INH(p[86])) ? `INH(p[86]) : y[83];
        y[84] = `C255;
        y[84] = (y[84] > `INH(p[12])) ? `INH(p[12]) : y[84];
        y[84] = (y[84] > `INH(p[85])) ? `INH(p[85]) : y[84];
        y[84] = (y[84] > p[86]) ? p[86] : y[84];
        y[85] = `C255;
        y[85] = (y[85] > `INH(p[84])) ? `INH(p[84]) : y[85];
        y[85] = (y[85] > `INH(p[86])) ? `INH(p[86]) : y[85];
        y[85] = (y[85] > p[87]) ? p[87] : y[85];
        y[86] = `C255;
        y[86] = (y[86] > `INH(p[2])) ? `INH(p[2]) : y[86];
        y[86] = (y[86] > p[81]) ? p[81] : y[86];
        y[86] = (y[86] > p[85]) ? p[85] : y[86];
        y[87] = `C255;
        y[87] = (y[87] > p[67]) ? p[67] : y[87];
        y[87] = (y[87] > `INH(p[83])) ? `INH(p[83]) : y[87];
        y[87] = (y[87] > `INH(p[87])) ? `INH(p[87]) : y[87];
        y[88] = `C255;
        y[88] = (y[88] > p[68]) ? p[68] : y[88];
        y[88] = (y[88] > `INH(p[88])) ? `INH(p[88]) : y[88];
        y[89] = `C255;
        y[89] = (y[89] > p[13]) ? p[13] : y[89];
        y[89] = (y[89] > `INH(p[69])) ? `INH(p[69]) : y[89];
        y[90] = `C255;
        y[90] = (y[90] > `INH(p[13])) ? `INH(p[13]) : y[90];
        y[90] = (y[90] > `INH(p[69])) ? `INH(p[69]) : y[90];
        y[90] = (y[90] > p[88]) ? p[88] : y[90];
        y[91] = `C255;
        y[91] = (y[91] > p[3]) ? p[3] : y[91];
        y[91] = (y[91] > `INH(p[68])) ? `INH(p[68]) : y[91];
        y[91] = (y[91] > `INH(p[88])) ? `INH(p[88]) : y[91];
        y[92] = `C255;
        y[92] = (y[92] > p[90]) ? p[90] : y[92];
        y[92] = (y[92] > `INH(p[92])) ? `INH(p[92]) : y[92];
        y[93] = `C255;
        y[93] = (y[93] > `INH(p[89])) ? `INH(p[89]) : y[93];
        y[93] = (y[93] > `INH(p[90])) ? `INH(p[90]) : y[93];
        y[93] = (y[93] > `INH(p[92])) ? `INH(p[92]) : y[93];
        y[93] = (y[93] > p[93]) ? p[93] : y[93];
        y[94] = `C255;
        y[94] = (y[94] > p[10]) ? p[10] : y[94];
        y[94] = (y[94] > `INH(p[95])) ? `INH(p[95]) : y[94];
        y[95] = `C255;
        y[95] = (y[95] > p[94]) ? p[94] : y[95];
        y[95] = (y[95] > `INH(p[96])) ? `INH(p[96]) : y[95];
        y[96] = `C255;
        y[96] = (y[96] > `INH(p[10])) ? `INH(p[10]) : y[96];
        y[96] = (y[96] > `INH(p[95])) ? `INH(p[95]) : y[96];
        y[96] = (y[96] > p[96]) ? p[96] : y[96];
        y[97] = `C255;
        y[97] = (y[97] > `INH(p[94])) ? `INH(p[94]) : y[97];
        y[97] = (y[97] > `INH(p[96])) ? `INH(p[96]) : y[97];
        y[97] = (y[97] > p[97]) ? p[97] : y[97];
        y[98] = `C255;
        y[98] = (y[98] > p[13]) ? p[13] : y[98];
        y[98] = (y[98] > `INH(p[99])) ? `INH(p[99]) : y[98];
        y[99] = `C255;
        y[99] = (y[99] > p[98]) ? p[98] : y[99];
        y[99] = (y[99] > `INH(p[100])) ? `INH(p[100]) : y[99];
        y[100] = `C255;
        y[100] = (y[100] > `INH(p[13])) ? `INH(p[13]) : y[100];
        y[100] = (y[100] > `INH(p[99])) ? `INH(p[99]) : y[100];
        y[100] = (y[100] > p[100]) ? p[100] : y[100];
        y[101] = `C255;
        y[101] = (y[101] > `INH(p[98])) ? `INH(p[98]) : y[101];
        y[101] = (y[101] > `INH(p[100])) ? `INH(p[100]) : y[101];
        y[101] = (y[101] > p[101]) ? p[101] : y[101];
        y[102] = `C255;
        y[102] = (y[102] > `INH(p[3])) ? `INH(p[3]) : y[102];
        y[102] = (y[102] > p[95]) ? p[95] : y[102];
        y[102] = (y[102] > p[99]) ? p[99] : y[102];
        y[103] = `C255;
        y[103] = (y[103] > p[92]) ? p[92] : y[103];
        y[103] = (y[103] > `INH(p[97])) ? `INH(p[97]) : y[103];
        y[103] = (y[103] > `INH(p[101])) ? `INH(p[101]) : y[103];
        y[104] = `C255;
        y[104] = (y[104] > p[91]) ? p[91] : y[104];
        y[104] = (y[104] > `INH(p[102])) ? `INH(p[102]) : y[104];
        y[105] = `C255;
        y[105] = (y[105] > p[14]) ? p[14] : y[105];
        y[105] = (y[105] > `INH(p[93])) ? `INH(p[93]) : y[105];
        y[106] = `C255;
        y[106] = (y[106] > `INH(p[14])) ? `INH(p[14]) : y[106];
        y[106] = (y[106] > `INH(p[93])) ? `INH(p[93]) : y[106];
        y[106] = (y[106] > p[102]) ? p[102] : y[106];
        y[107] = `C255;
        y[107] = (y[107] > p[4]) ? p[4] : y[107];
        y[107] = (y[107] > `INH(p[91])) ? `INH(p[91]) : y[107];
        y[107] = (y[107] > `INH(p[102])) ? `INH(p[102]) : y[107];
        y[108] = `C255;
        y[108] = (y[108] > p[104]) ? p[104] : y[108];
        y[108] = (y[108] > `INH(p[106])) ? `INH(p[106]) : y[108];
        y[109] = `C255;
        y[109] = (y[109] > `INH(p[103])) ? `INH(p[103]) : y[109];
        y[109] = (y[109] > `INH(p[104])) ? `INH(p[104]) : y[109];
        y[109] = (y[109] > `INH(p[106])) ? `INH(p[106]) : y[109];
        y[109] = (y[109] > p[107]) ? p[107] : y[109];
        y[110] = `C255;
        y[110] = (y[110] > p[14]) ? p[14] : y[110];
        y[110] = (y[110] > `INH(p[109])) ? `INH(p[109]) : y[110];
        y[111] = `C255;
        y[111] = (y[111] > p[108]) ? p[108] : y[111];
        y[111] = (y[111] > `INH(p[110])) ? `INH(p[110]) : y[111];
        y[112] = `C255;
        y[112] = (y[112] > `INH(p[14])) ? `INH(p[14]) : y[112];
        y[112] = (y[112] > `INH(p[109])) ? `INH(p[109]) : y[112];
        y[112] = (y[112] > p[110]) ? p[110] : y[112];
        y[113] = `C255;
        y[113] = (y[113] > `INH(p[108])) ? `INH(p[108]) : y[113];
        y[113] = (y[113] > `INH(p[110])) ? `INH(p[110]) : y[113];
        y[113] = (y[113] > p[111]) ? p[111] : y[113];
        y[114] = `C255;
        y[114] = (y[114] > p[15]) ? p[15] : y[114];
        y[114] = (y[114] > `INH(p[113])) ? `INH(p[113]) : y[114];
        y[115] = `C255;
        y[115] = (y[115] > p[112]) ? p[112] : y[115];
        y[115] = (y[115] > `INH(p[114])) ? `INH(p[114]) : y[115];
        y[116] = `C255;
        y[116] = (y[116] > `INH(p[15])) ? `INH(p[15]) : y[116];
        y[116] = (y[116] > `INH(p[113])) ? `INH(p[113]) : y[116];
        y[116] = (y[116] > p[114]) ? p[114] : y[116];
        y[117] = `C255;
        y[117] = (y[117] > `INH(p[112])) ? `INH(p[112]) : y[117];
        y[117] = (y[117] > `INH(p[114])) ? `INH(p[114]) : y[117];
        y[117] = (y[117] > p[115]) ? p[115] : y[117];
        y[118] = `C255;
        y[118] = (y[118] > `INH(p[4])) ? `INH(p[4]) : y[118];
        y[118] = (y[118] > p[109]) ? p[109] : y[118];
        y[118] = (y[118] > p[113]) ? p[113] : y[118];
        y[119] = `C255;
        y[119] = (y[119] > p[106]) ? p[106] : y[119];
        y[119] = (y[119] > `INH(p[111])) ? `INH(p[111]) : y[119];
        y[119] = (y[119] > `INH(p[115])) ? `INH(p[115]) : y[119];
        y[120] = `C255;
        y[120] = (y[120] > p[105]) ? p[105] : y[120];
        y[120] = (y[120] > `INH(p[116])) ? `INH(p[116]) : y[120];
        y[121] = `C255;
        y[121] = (y[121] > p[16]) ? p[16] : y[121];
        y[121] = (y[121] > `INH(p[107])) ? `INH(p[107]) : y[121];
        y[122] = `C255;
        y[122] = (y[122] > `INH(p[16])) ? `INH(p[16]) : y[122];
        y[122] = (y[122] > `INH(p[107])) ? `INH(p[107]) : y[122];
        y[122] = (y[122] > p[116]) ? p[116] : y[122];
        y[123] = `C255;
        y[123] = (y[123] > p[5]) ? p[5] : y[123];
        y[123] = (y[123] > `INH(p[105])) ? `INH(p[105]) : y[123];
        y[123] = (y[123] > `INH(p[116])) ? `INH(p[116]) : y[123];


		if(y[5]>`C0)
                y[0] = `C0;
        if(y[6]>`C0)
                y[7] = `C0;
        if(y[8]>`C0)
                y[9] = `C0;
        if(y[10]>`C0)
                y[11] = `C0;
        if(y[12]>`C0)
                y[14] = `C0;
        if(y[13]>`C0)
                y[14] = `C0;
        if(y[15]>`C0)
                y[16] = `C0;
        if(y[17]>`C0)
                y[18] = `C0;
        if(y[17]>`C0)
                y[19] = `C0;
        if(y[34]>`C0)
                y[1] = `C0;
        if(y[35]>`C0)
                y[36] = `C0;
        if(y[37]>`C0)
                y[38] = `C0;
        if(y[39]>`C0)
                y[40] = `C0;
        if(y[41]>`C0)
                y[43] = `C0;
        if(y[42]>`C0)
                y[43] = `C0;
        if(y[44]>`C0)
                y[45] = `C0;
        if(y[46]>`C0)
                y[47] = `C0;
        if(y[46]>`C0)
                y[48] = `C0;
        if(y[63]>`C0)
                y[2] = `C0;
        if(y[64]>`C0)
                y[65] = `C0;
        if(y[66]>`C0)
                y[67] = `C0;
        if(y[68]>`C0)
                y[69] = `C0;
        if(y[70]>`C0)
                y[72] = `C0;
        if(y[71]>`C0)
                y[72] = `C0;
        if(y[73]>`C0)
                y[74] = `C0;
        if(y[75]>`C0)
                y[76] = `C0;
        if(y[75]>`C0)
                y[77] = `C0;


                if(y[0]>`C0) begin
                        p[22] = p[22] - y[0];
                        p[19] = p[19] + y[0];
                end else 
                if(y[1]>`C0) begin
                        p[46] = p[46] - y[1];
                        p[43] = p[43] + y[1];
                end else
  // required to process
                if(y[2]>`C0) begin
                        p[70] = p[70] - y[2];
                        p[67] = p[67] + y[2];
                end else
                if(y[3]>`C0) begin
                        p[89] = p[89] - y[3];
                        p[91] = p[91] + y[3];
                end else
                if(y[4]>`C0) begin
                        p[103] = p[103] - y[4];
                        p[105] = p[105] + y[4];
                end else
                if(y[5]>`C0) begin
                        p[23] = p[23] - y[5];
                        p[19] = p[19] + y[5];
                end else
                if(y[6]>`C0) begin
                        p[17] = p[17] - y[6];
                end else
                if(y[7]>`C0) begin
                        p[21] = p[21] - y[7];
                        p[23] = p[23] + y[7];
                end else
                if(y[8]>`C0) begin
                        p[18] = p[18] - y[8]*`C2;
                        p[24] = p[24] + y[8];
                end else
                if(y[9]>`C0) begin
                        p[25] = p[25] - y[9];
                        p[22] = p[22] + y[9];
                end else
                if(y[10]>`C0) begin
                        p[18] = p[18] - y[10];
                        p[27] = p[27] - y[10];
                        p[26] = p[26] + y[10];
                end else
                if(y[11]>`C0) begin
                        p[28] = p[28] - y[11];
                        p[25] = p[25] + y[11];
                end else
                if(y[12]>`C0) begin
                        p[17] = p[17] - y[12];
                        p[20] = p[20] + y[12];
                        p[29] = p[29] + y[12];
                end else
                if(y[13]>`C0) begin
                        p[17] = p[17] - y[13];
                        p[29] = p[29] + y[13];
                end else
                if(y[14]>`C0) begin
                        p[30] = p[30] - y[14];
                        p[28] = p[28] + y[14];
                end else
                if(y[15]>`C0) begin
                        p[24] = p[24] - y[15];
                        p[18] = p[18] + y[15];
                end else
                if(y[16]>`C0) begin
                        p[31] = p[31] - y[16];
                        p[30] = p[30] + y[16];
                end else
                if(y[17]>`C0) begin
                        p[29] = p[29] - y[17];
                        p[17] = p[17] + y[17]*`C2;
                end else
                if(y[18]>`C0) begin
                        p[19] = p[19] - y[18];
                        p[26] = p[26] - y[18];
                        p[27] = p[27] + y[18];
                        p[31] = p[31] + y[18];
                end else
                if(y[19]>`C0) begin
                        p[19] = p[19] - y[19];
                        p[31] = p[31] + y[19];
                end else
                if(y[20]>`C0) begin
                        p[6] = p[6] - y[20];
                        p[17] = p[17] + y[20];
                        p[32] = p[32] + y[20];
                end else
                if(y[21]>`C0) begin
                        p[32] = p[32] - y[21];
                        p[6] = p[6] + y[21];
                end else
                if(y[22]>`C0) begin
                        
                        p[34] = p[34] - y[22];
                        p[33] = p[33] + y[22];
                end else
                if(y[23]>`C0) begin
                        
                        p[35] = p[35] - y[23];
                        p[34] = p[34] + y[23];
                end else
                if(y[24]>`C0) begin
//                        y[] = y[24];
                        p[7] = p[7] - y[24];
                        p[18] = p[18] + y[24];
                        p[36] = p[36] + y[24];
                end else
                if(y[25]>`C0) begin
//                        y[] = y[25];
                        p[36] = p[36] - y[25];
                        p[7] = p[7] + y[25];
                end else
                if(y[26]>`C0) begin
//                        y[] = y[26];
                        p[38] = p[38] - y[26];
                        p[37] = p[37] + y[26];
                end else
                if(y[27]>`C0) begin
//                        y[] = y[27];
                        p[39] = p[39] - y[27];
                        p[38] = p[38] + y[27];
                end else
                if(y[28]>`C0) begin
//                        y[] = y[28];
                        p[33] = p[33] - y[28];
                        p[37] = p[37] - y[28];
                        p[0] = p[0] + y[28];
                end else
                if(y[29]>`C0) begin
//                        y[] = y[29];
                        p[19] = p[19] - y[29];
                        p[35] = p[35] + y[29];
                        p[39] = p[39] + y[29];
                end else
                if(y[30]>`C0) begin
//                        y[] = y[30];
                        p[20] = p[20] - y[30];
                        p[8] = p[8] + y[30];
                end else
                if(y[31]>`C0) begin
//                        y[] = y[31];
                        p[8] = p[8] - y[31];
                end else
                if(y[32]>`C0) begin
//                        y[] = y[32];
                        p[40] = p[40] - y[32];
                        p[21] = p[21] + y[32];
                end else
                if(y[33]>`C0) begin
//                        y[] = y[33];
                        p[1] = p[1] - y[33];
                        p[40] = p[40] + y[33];
                end else
                if(y[34]>`C0) begin
//                        y[] = y[34];
                        p[47] = p[47] - y[34];
                        p[43] = p[43] + y[34];
                end else
                if(y[35]>`C0) begin
//                        y[] = y[35];
                        p[41] = p[41] - y[35];
                end else
                if(y[36]>`C0) begin
//                        y[] = y[36];
                        p[45] = p[45] - y[36];
                        p[47] = p[47] + y[36];
                end else
                if(y[37]>`C0) begin
//                        y[] = y[37];
                        p[42] = p[42] - y[37]*`C2;
                        p[48] = p[48] + y[37];
                end else
                if(y[38]>`C0) begin
//                        y[] = y[38];
                        p[49] = p[49] - y[38];
                        p[46] = p[46] + y[38];
                end else
                if(y[39]>`C0) begin
//                        y[] = y[39];
                        p[42] = p[42] - y[39];
                        p[51] = p[51] - y[39];
                        p[50] = p[50] + y[39];
                end else
                if(y[40]>`C0) begin
//                        y[] = y[40];
                        p[52] = p[52] - y[40];
                        p[49] = p[49] + y[40];
                end else
                if(y[41]>`C0) begin
//                        y[] = y[41];
                        p[41] = p[41] - y[41];
                        p[44] = p[44] + y[41];
                        p[53] = p[53] + y[41];
                end else
                if(y[42]>`C0) begin
//                        y[] = y[42];
                        p[41] = p[41] - y[42];
                        p[53] = p[53] + y[42];
                end else
                if(y[43]>`C0) begin
//                        y[] = y[43];
                        p[54] = p[54] - y[43];
                        p[52] = p[52] + y[43];
                end else
                if(y[44]>`C0) begin
//                        y[] = y[44];
                        p[48] = p[48] - y[44];
                        p[42] = p[42] + y[44];
                end else
                if(y[45]>`C0) begin
//                        y[] = y[45];
                        p[55] = p[55] - y[45];
                        p[54] = p[54] + y[45];
                end else
                if(y[46]>`C0) begin
//                        y[] = y[46];
                        p[53] = p[53] - y[46];
                        p[41] = p[41] + y[46]*`C2;
                end else
                if(y[47]>`C0) begin
//                        y[] = y[47];
                        p[43] = p[43] - y[47];
                        p[50] = p[50] - y[47];
                        p[51] = p[51] + y[47];
                        p[55] = p[55] + y[47];
                end else
                if(y[48]>`C0) begin
//                        y[] = y[48];
                        p[43] = p[43] - y[48];
                        p[55] = p[55] + y[48];
                end else
                if(y[49]>`C0) begin
//                        y[] = y[49];
                        p[8] = p[8] - y[49];
                        p[41] = p[41] + y[49];
                        p[56] = p[56] + y[49];
                end else
                if(y[50]>`C0) begin
//                        y[] = y[50];
                        p[56] = p[56] - y[50];
                        p[8] = p[8] + y[50];
                end else
                if(y[51]>`C0) begin
//                        y[] = y[51];
                        p[58] = p[58] - y[51];
                        p[57] = p[57] + y[51];
                end else
                if(y[52]>`C0) begin
//                        y[] = y[52];
                        p[59] = p[59] - y[52];
                        p[58] = p[58] + y[52];
                end else
                if(y[53]>`C0) begin
//                        y[] = y[53];
                        p[9] = p[9] - y[53];
                        p[42] = p[42] + y[53];
                        p[60] = p[60] + y[53];
                end else
                if(y[54]>`C0) begin
//                        y[] = y[54];
                        p[60] = p[60] - y[54];
                        p[9] = p[9] + y[54];
                end else
                if(y[55]>`C0) begin
//                        y[] = y[55];
                        p[62] = p[62] - y[55];
                        p[61] = p[61] + y[5];
                end else
                if(y[56]>`C0) begin
//                        y[] = y[56];
                        p[63] = p[63] - y[56];
                        p[62] = p[62] + y[56];
                end else
                if(y[57]>`C0) begin
//                        y[] = y[57];
                        p[57] = p[57] - y[57];
                        p[61] = p[61] - y[57];
                        p[1] = p[1] + y[57];
                end else
                if(y[58]>`C0) begin
//                        y[] = y[58];
                        p[43] = p[43] - y[58];
                        p[59] = p[59] + y[58];
                        p[63] = p[63] + y[58];
                end else
                if(y[59]>`C0) begin
//                        y[] = y[59];
                        p[44] = p[44] - y[59];
                        p[10] = p[10] + y[59];
                end else
                if(y[60]>`C0) begin
//                        y[] = y[60];
                        p[10] = p[10] - y[60];
                end else
                if(y[61]>`C0) begin
//                        y[] = y[61];
                        p[64] = p[64] - y[61];
                        p[45] = p[45] + y[61];
                end else
                if(y[62]>`C0) begin
//                        y[] = y[62];
                        p[2] = p[2] - y[62];
                        p[64] = p[64] + y[62];
                end else
                if(y[63]>`C0) begin
//                        y[] = y[63];
                        p[71] = p[71] - y[63];
                        p[67] = p[67] + y[63];
                end else
                if(y[64]>`C0) begin
//                        y[] = y[64];
                        p[65] = p[65] - y[64];
                end else
                if(y[65]>`C0) begin
//                        y[] = y[65];
                        p[69] = p[69] - y[65];
                        p[71] = p[71] + y[65];
                end else
                if(y[66]>`C0) begin
//                        y[] = y[66];
                        p[66] = p[66] - y[66]*`C2;
                        p[72] = p[72] + y[66];
                end else
                if(y[67]>`C0) begin
//                        y[] = y[67];
                        p[73] = p[73] - y[67];
                        p[70] = p[70] + y[67];
                end else
                if(y[68]>`C0) begin
//                        y[] = y[68];
                        p[66] = p[66] - y[68];
                        p[75] = p[75] - y[68];
                        p[74] = p[74] + y[68];
                end else
                if(y[69]>`C0) begin
//                        y[] = y[69];
                        p[76] = p[76] - y[69];
                        p[73] = p[73] + y[69];
                end else
                if(y[70]>`C0) begin
//                        y[] = y[70];
                        p[65] = p[65] - y[70];
                        p[68] = p[68] + y[70];
                        p[77] = p[77] + y[70];
                end else
                if(y[71]>`C0) begin
//                        y[] = y[71];
                        p[65] = p[65] - y[71];
                        p[77] = p[77] + y[71];
                end else
                if(y[72]>`C0) begin
//                        y[] = y[72];
                        p[78] = p[78] - y[72];
                        p[76] = p[76] + y[72];
                end else
                if(y[73]>`C0) begin
//                        y[] = y[73];
                        p[72] = p[72] - y[73];
                        p[66] = p[66] + y[73];
                end else
                if(y[74]>`C0) begin
//                        y[] = y[74];
                        p[79] = p[79] - y[74];
                        p[78] = p[78] + y[74];
                end else
                if(y[75]>`C0) begin
//                        y[] = y[75];
                        p[77] = p[77] - y[75];
                        p[65] = p[65] + y[75]*`C2;
                end else
                if(y[76]>`C0) begin
//                        y[] = y[76];
                        p[67] = p[67] - y[76];
                        p[74] = p[74] - y[76];
                        p[75] = p[75] + y[76];
                        p[79] = p[79] + y[76];
                end else
                if(y[77]>`C0) begin
//                        y[] = y[77];
                        p[67] = p[67] - y[77];
                        p[79] = p[79] + y[77];
                end else
                if(y[78]>`C0) begin
//                        y[] = y[78];
                        p[11] = p[11] - y[78];
                        p[65] = p[65] + y[78];
                        p[80] = p[80] + y[78];
                end else
                if(y[79]>`C0) begin
//                        y[] = y[79];
                        p[80] = p[80] - y[79];
                        p[11] = p[11] + y[79];
                end else
                if(y[80]>`C0) begin
//                        y[] = y[80];
                        p[82] = p[82] - y[80];
                        p[81] = p[81] + y[80];
                end else
                if(y[81]>`C0) begin
//                        y[] = y[81];
                        p[83] = p[83] - y[81];
                        p[82] = p[82] + y[81];
                end else
                if(y[82]>`C0) begin
//                        y[] = y[82];
                        p[12] = p[12] - y[82];
                        p[66] = p[66] + y[82];
                        p[84] = p[84] + y[82];
                end else
                if(y[83]>`C0) begin
//                        y[] = y[83];
                        p[84] = p[84] - y[83];
                        p[12] = p[12] + y[83];
                end else
                if(y[84]>`C0) begin
//                        y[] = y[84];
                        p[86] = p[86] - y[84];
                        p[85] = p[85] + y[84];
                end else
                if(y[85]>`C0) begin
//                        y[] = y[85];
                        p[87] = p[87] - y[85];
                        p[86] = p[86] + y[85];
                end else
                if(y[86]>`C0) begin
//                        y[] = y[86];
                        p[81] = p[81] - y[86];
                        p[85] = p[85] - y[86];
                        p[2] = p[2] + y[86];
                end else
                if(y[87]>`C0) begin
//                        y[] = y[87];
                        p[67] = p[67] - y[87];
                        p[83] = p[83] + y[87];
                        p[87] = p[87] + y[87];
                end else
                if(y[88]>`C0) begin
//                        y[] = y[88];
                        p[68] = p[68] - y[88];
                        p[13] = p[13] + y[88];
                end else
                if(y[89]>`C0) begin
//                        y[] = y[89];
                        p[13] = p[13] - y[89];
                end else
                if(y[90]>`C0) begin
//                        y[] = y[90];
                        p[88] = p[88] - y[90];
                        p[69] = p[69] + y[90];
                end else
                if(y[91]>`C0) begin
//                        y[] = y[91];
                        p[3] = p[3] - y[91];
                        p[88] = p[88] + y[91];
                end else
                if(y[92]>`C0) begin
//                        y[] = y[92];
                        p[90] = p[90] - y[92];
                        p[91] = p[91] + y[92];
                end else
                if(y[93]>`C0) begin
//                        y[] = y[93];
                        p[93] = p[93] - y[93];
                        p[92] = p[92] + y[93];
                end else
                if(y[94]>`C0) begin
//                        y[] = y[94];
                        p[10] = p[10] - y[94];
                        p[89] = p[89] + y[94];
                        p[94] = p[94] + y[94];
                end else
                if(y[95]>`C0) begin
//                        y[] = y[95];
                        p[94] = p[94] - y[95];
                        p[10] = p[10] + y[95];
                end else
                if(y[96]>`C0) begin
//                        y[] = y[96];
                        p[96] = p[96] - y[96];
                        p[95] = p[95] + y[96];
                end else
                if(y[97]>`C0) begin
//                        y[] = y[97];
                        p[97] = p[97] - y[97];
                        p[96] = p[96] + y[97];
                end else
                if(y[98]>`C0) begin
//                        y[] = y[98];
                        p[13] = p[13] - y[98];
                        p[90] = p[90] + y[98];
                        p[98] = p[98] + y[98];
                end else
                if(y[99]>`C0) begin
//                        y[] = y[99];
                        p[98] = p[98] - y[99];
                        p[13] = p[13] + y[99];
                end else
                if(y[100]>`C0) begin
//                        y[] = y[100];
                        p[100] = p[100] - y[100];
                        p[99] = p[99] + y[100];
                end else
                if(y[101]>`C0) begin
//                        y[] = y[101];
                        p[101] = p[101] - y[101];
                        p[100] = p[100] + y[101];
                end else
                if(y[102]>`C0) begin
//                        y[] = y[102];
                        p[95] = p[95] - y[102];
                        p[99] = p[99] - y[102];
                        p[3] = p[3] + y[102];
                end else
                if(y[103]>`C0) begin
//                        y[] = y[103];
                        p[92] = p[92] - y[103];
                        p[97] = p[97] + y[103];
                        p[101] = p[101] + y[103];
                end else
                if(y[104]>`C0) begin
//                        y[] = y[104];
                        p[91] = p[91] - y[104];
                        p[14] = p[14] + y[104];
                end else
                if(y[105]>`C0) begin
//                        y[] = y[105];
                        p[14] = p[14] - y[105];
                end else
                if(y[106]>`C0) begin
//                        y[] = y[106];
                        p[102] = p[102] - y[106];
                        p[93] = p[93] + y[106];
                end else
                if(y[107]>`C0) begin
//                        y[] = y[107];
                        p[4] = p[4] - y[107];
                        p[102] = p[102] + y[107];
                end else
                if(y[108]>`C0) begin
//                        y[] = y[108];
                        p[104] = p[104] - y[108];
                        p[105] = p[105] + y[108];
                end else
                if(y[109]>`C0) begin
                        p[107] = p[107] - y[109];
                        p[106] = p[106] + y[109];
                end else
                if(y[110]>`C0) begin
                        p[14] = p[14] - y[110];
                        p[103] = p[103] + y[110];
                        p[108] = p[108] + y[110];
                end else
                if(y[111]>`C0) begin
                        p[108] = p[108] - y[111];
                        p[14] = p[14] + y[111];
                end else
                if(y[112]>`C0) begin
                        p[110] = p[110] - y[112];
                        p[109] = p[109] + y[112];
                end else
                if(y[113]>`C0) begin
                        p[111] = p[111] - y[113];
                        p[110] = p[110] + y[113];
                end else
                if(y[114]>`C0) begin
                        p[15] = p[15] - y[114];
                        p[104] = p[104] + y[114];
                        p[112] = p[112] + y[114];
                end else
                if(y[115]>`C0) begin
                        p[112] = p[112] - y[115];
                        p[15] = p[15] + y[115];
                end else
                if(y[116]>`C0) begin
                        p[114] = p[114] - y[116];
                        p[113] = p[113] + y[116];
                end else
                if(y[117]>`C0) begin
                        p[115] = p[115] - y[117];
                        p[114] = p[114] + y[117];
                end else
                if(y[118]>`C0) begin
                        p[109] = p[109] - y[118];
                        p[113] = p[113] - y[118];
                        p[4] = p[4] + y[118];
                end else
                if(y[119]>`C0) begin
                        p[106] = p[106] - y[119];
                        p[111] = p[111] + y[119];
                        p[115] = p[115] + y[119];
                end else
                if(y[120]>`C0) begin
                        p[105] = p[105] - y[120];
                        p[16] = p[16] + y[120];
                end else
                if(y[121]>`C0) begin
                        p[16] = p[16] - y[121];
                end else
                if(y[122]>`C0) begin
                        p[116] = p[116] - y[122];
                        p[107] = p[107] + y[122];
                end else
                if(y[123]>`C0) begin
                        p[5] = p[5] - y[123];
                        p[116] = p[116] + y[123];
                end

  // end required to process
        

//        if(tf!=`C0) begin 
//            led = 6'b000000; 
//        end else begin 
            led = ~(p[16][5:0]); 
//        end
        
end

endmodule
