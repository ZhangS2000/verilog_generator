module sn(
        input clk,
        output reg [5:0] led
);
`define INH(place) ((place) == 0 ? 4095 : 0)
reg [10:0] p[670:0]={0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,8,2,0,2,0,2,0,2,0,2,0,2,0,5,2,0,2,0,2,0,2,0,2,0,0,1,2,0,2,0,2,0,2,0,0,10,2,0,2,0,2,0,0,5,2,0,2,0,0,9,2,0,0,9,0,0,0,1,0,1,1,1,0,1,0,1,1,0,1,1,0,1,1,1,0,1,1,1,1,0,0,1,0,1,1,1,0,1,0,1,1,0,1,1,0,1,1,1,0,1,1,1,1,0,0,1,0,1,1,1,0,1,0,1,1,0,1,1,0,1,1,1,0,1,1,1,1,0,0,1,0,1,1,1,0,1,0,1,1,0,1,1,0,1,1,1,0,1,1,1,1,0,0,1,0,1,1,1,0,1,0,1,1,0,1,1,0,1,1,1,0,1,1,1,1,0,0,1,0,1,1,1,0,1,0,1,1,0,1,1,0,1,1,1,0,1,1,1,1,0,0,1,0,1,1,1,0,1,0,1,1,0,1,1,0,1,1,1,0,1,1,1,1,0,0,1,0,1,1,1,0,1,0,1,1,0,1,1,0,1,1,1,0,1,1,1,1,0,0,1,0,1,1,1,0,1,0,1,1,0,1,1,0,1,1,1,0,1,1,1,1,0,0,1,0,1,1,1,0,1,0,1,1,0,1,1,0,1,1,1,0,1,1,1,1,0,0,1,0,1,1,1,0,1,0,1,1,0,1,1,0,1,1,1,0,1,1,1,1,0,0,0,1,1,0,1,1,1,0,1,1,1,1,0,0,1,0,1,1,1,0,1,0,1,1,0,1,1,0,1,1,1,0,1,1,1,1,0,0,1,0,1,1,1,0,1,0,1,1,0,1,1,0,1,1,1,0,1,1,1,1,0,0,1,0,1,1,1,0,1,0,1,1,0,1,1,0,1,1,1,0,1,1,1,1,0,0,1,0,1,1,1,0,1,0,1,1,0,1,1,0,1,1,1,0,1,1,1,1,0,0,0,1,1,0,1,1,1,0,1,1,1,1,0,0,1,0,1,1,1,0,1,0,1,1,0,1,1,0,1,1,1,0,1,1,1,1,0,0,1,0,1,1,1,0,1,0,1,1,0,1,1,0,1,1,1,0,1,1,1,1,0,0,1,0,1,1,1,0,1,0,1,1,0,1,1,0,1,1,1,0,1,1,1,1,0,0,0,1,1,0,1,1,1,0,1,1,1,1,0,0,1,0,1,1,1,0,1,0,1,1,0,1,1,0,1,1,1,0,1,1,1,1,0,0,1,0,1,1,1,0,1,0,1,1,0,1,1,0,1,1,1,0,1,1,1,1,0,0,0,1,1,0,1,1,1,0,1,1,1,1,0,0,1,0,1,1,1,0,1,0,1,1,0,1,1,0,1,1,1,0,1,1,1,1,0,0,0,1,1,0,1,1,1,0,1,1,1,1,0,0,0,1,1,0,1,1,1,0,1,1,1,1};
reg [10:0] f[731:0];
reg [10:0] tf;
reg [10:0] tc;
always @(posedge clk) begin
        f[0] = 4095;
        f[0] = (f[0] >= `INH(p[85])) ? `INH(p[85]) : f[0];
        f[0] = (f[0] > p[88]) ? p[88] : f[0];
        f[1] = 4095;
        f[1] = (f[1] >= `INH(p[109])) ? `INH(p[109]) : f[1];
        f[1] = (f[1] > p[112]) ? p[112] : f[1];
        f[2] = 4095;
        f[2] = (f[2] >= `INH(p[133])) ? `INH(p[133]) : f[2];
        f[2] = (f[2] > p[136]) ? p[136] : f[2];
        f[3] = 4095;
        f[3] = (f[3] >= `INH(p[157])) ? `INH(p[157]) : f[3];
        f[3] = (f[3] > p[160]) ? p[160] : f[3];
        f[4] = 4095;
        f[4] = (f[4] >= `INH(p[181])) ? `INH(p[181]) : f[4];
        f[4] = (f[4] > p[184]) ? p[184] : f[4];
        f[5] = 4095;
        f[5] = (f[5] >= `INH(p[205])) ? `INH(p[205]) : f[5];
        f[5] = (f[5] > p[208]) ? p[208] : f[5];
        f[6] = 4095;
        f[6] = (f[6] >= `INH(p[229])) ? `INH(p[229]) : f[6];
        f[6] = (f[6] > p[232]) ? p[232] : f[6];
        f[7] = 4095;
        f[7] = (f[7] >= `INH(p[253])) ? `INH(p[253]) : f[7];
        f[7] = (f[7] > p[256]) ? p[256] : f[7];
        f[8] = 4095;
        f[8] = (f[8] >= `INH(p[277])) ? `INH(p[277]) : f[8];
        f[8] = (f[8] > p[280]) ? p[280] : f[8];
        f[9] = 4095;
        f[9] = (f[9] >= `INH(p[301])) ? `INH(p[301]) : f[9];
        f[9] = (f[9] > p[304]) ? p[304] : f[9];
        f[10] = 4095;
        f[10] = (f[10] >= `INH(p[325])) ? `INH(p[325]) : f[10];
        f[10] = (f[10] > p[328]) ? p[328] : f[10];
        f[11] = 4095;
        f[11] = (f[11] > p[347]) ? p[347] : f[11];
        f[11] = (f[11] >= `INH(p[350])) ? `INH(p[350]) : f[11];
        f[12] = 4095;
        f[12] = (f[12] >= `INH(p[363])) ? `INH(p[363]) : f[12];
        f[12] = (f[12] > p[366]) ? p[366] : f[12];
        f[13] = 4095;
        f[13] = (f[13] >= `INH(p[387])) ? `INH(p[387]) : f[13];
        f[13] = (f[13] > p[390]) ? p[390] : f[13];
        f[14] = 4095;
        f[14] = (f[14] >= `INH(p[411])) ? `INH(p[411]) : f[14];
        f[14] = (f[14] > p[414]) ? p[414] : f[14];
        f[15] = 4095;
        f[15] = (f[15] >= `INH(p[435])) ? `INH(p[435]) : f[15];
        f[15] = (f[15] > p[438]) ? p[438] : f[15];
        f[16] = 4095;
        f[16] = (f[16] > p[457]) ? p[457] : f[16];
        f[16] = (f[16] >= `INH(p[460])) ? `INH(p[460]) : f[16];
        f[17] = 4095;
        f[17] = (f[17] >= `INH(p[473])) ? `INH(p[473]) : f[17];
        f[17] = (f[17] > p[476]) ? p[476] : f[17];
        f[18] = 4095;
        f[18] = (f[18] >= `INH(p[497])) ? `INH(p[497]) : f[18];
        f[18] = (f[18] > p[500]) ? p[500] : f[18];
        f[19] = 4095;
        f[19] = (f[19] >= `INH(p[521])) ? `INH(p[521]) : f[19];
        f[19] = (f[19] > p[524]) ? p[524] : f[19];
        f[20] = 4095;
        f[20] = (f[20] > p[543]) ? p[543] : f[20];
        f[20] = (f[20] >= `INH(p[546])) ? `INH(p[546]) : f[20];
        f[21] = 4095;
        f[21] = (f[21] >= `INH(p[559])) ? `INH(p[559]) : f[21];
        f[21] = (f[21] > p[562]) ? p[562] : f[21];
        f[22] = 4095;
        f[22] = (f[22] >= `INH(p[583])) ? `INH(p[583]) : f[22];
        f[22] = (f[22] > p[586]) ? p[586] : f[22];
        f[23] = 4095;
        f[23] = (f[23] > p[605]) ? p[605] : f[23];
        f[23] = (f[23] >= `INH(p[608])) ? `INH(p[608]) : f[23];
        f[24] = 4095;
        f[24] = (f[24] >= `INH(p[621])) ? `INH(p[621]) : f[24];
        f[24] = (f[24] > p[624]) ? p[624] : f[24];
        f[25] = 4095;
        f[25] = (f[25] > p[643]) ? p[643] : f[25];
        f[25] = (f[25] >= `INH(p[646])) ? `INH(p[646]) : f[25];
        f[26] = 4095;
        f[26] = (f[26] > p[657]) ? p[657] : f[26];
        f[26] = (f[26] >= `INH(p[660])) ? `INH(p[660]) : f[26];
        f[27] = 4095;
        f[27] = (f[27] >= `INH(p[84])) ? `INH(p[84]) : f[27];
        f[27] = (f[27] >= `INH(p[85])) ? `INH(p[85]) : f[27];
        f[27] = (f[27] > p[89]) ? p[89] : f[27];
        f[28] = 4095;
        f[28] = (f[28] > p[83]) ? p[83] : f[28];
        f[28] = (f[28] >= `INH(p[89])) ? `INH(p[89]) : f[28];
        f[29] = 4095;
        f[29] = (f[29] > p[87]) ? p[87] : f[29];
        f[29] = (f[29] >= `INH(p[89])) ? `INH(p[89]) : f[29];
        f[30] = 4095;
        f[30] = (f[30] >= p[84]/2) ? p[84]/2 : f[30];
        f[30] = (f[30] >= `INH(p[88])) ? `INH(p[88]) : f[30];
        f[31] = 4095;
        f[31] = (f[31] >= `INH(p[88])) ? `INH(p[88]) : f[31];
        f[31] = (f[31] > p[91]) ? p[91] : f[31];
        f[32] = 4095;
        f[32] = (f[32] > p[84]) ? p[84] : f[32];
        f[32] = (f[32] >= `INH(p[91])) ? `INH(p[91]) : f[32];
        f[32] = (f[32] > p[93]) ? p[93] : f[32];
        f[33] = 4095;
        f[33] = (f[33] >= `INH(p[91])) ? `INH(p[91]) : f[33];
        f[33] = (f[33] > p[94]) ? p[94] : f[33];
        f[34] = 4095;
        f[34] = (f[34] > p[83]) ? p[83] : f[34];
        f[34] = (f[34] >= `INH(p[93])) ? `INH(p[93]) : f[34];
        f[34] = (f[34] >= `INH(p[94])) ? `INH(p[94]) : f[34];
        f[35] = 4095;
        f[35] = (f[35] > p[83]) ? p[83] : f[35];
        f[35] = (f[35] >= `INH(p[92])) ? `INH(p[92]) : f[35];
        f[35] = (f[35] >= `INH(p[94])) ? `INH(p[94]) : f[35];
        f[36] = 4095;
        f[36] = (f[36] >= `INH(p[94])) ? `INH(p[94]) : f[36];
        f[36] = (f[36] > p[96]) ? p[96] : f[36];
        f[37] = 4095;
        f[37] = (f[37] > p[90]) ? p[90] : f[37];
        f[37] = (f[37] >= `INH(p[96])) ? `INH(p[96]) : f[37];
        f[38] = 4095;
        f[38] = (f[38] >= `INH(p[96])) ? `INH(p[96]) : f[38];
        f[38] = (f[38] > p[97]) ? p[97] : f[38];
        f[39] = 4095;
        f[39] = (f[39] > p[95]) ? p[95] : f[39];
        f[39] = (f[39] >= `INH(p[97])) ? `INH(p[97]) : f[39];
        f[40] = 4095;
        f[40] = (f[40] > p[85]) ? p[85] : f[40];
        f[40] = (f[40] > p[92]) ? p[92] : f[40];
        f[40] = (f[40] >= `INH(p[93])) ? `INH(p[93]) : f[40];
        f[40] = (f[40] >= `INH(p[97])) ? `INH(p[97]) : f[40];
        f[41] = 4095;
        f[41] = (f[41] > p[85]) ? p[85] : f[41];
        f[41] = (f[41] >= `INH(p[92])) ? `INH(p[92]) : f[41];
        f[41] = (f[41] >= `INH(p[97])) ? `INH(p[97]) : f[41];
        f[42] = 4095;
        f[42] = (f[42] > p[28]) ? p[28] : f[42];
        f[42] = (f[42] >= `INH(p[99])) ? `INH(p[99]) : f[42];
        f[43] = 4095;
        f[43] = (f[43] > p[98]) ? p[98] : f[43];
        f[43] = (f[43] >= `INH(p[100])) ? `INH(p[100]) : f[43];
        f[44] = 4095;
        f[44] = (f[44] >= `INH(p[28])) ? `INH(p[28]) : f[44];
        f[44] = (f[44] >= `INH(p[99])) ? `INH(p[99]) : f[44];
        f[44] = (f[44] > p[100]) ? p[100] : f[44];
        f[45] = 4095;
        f[45] = (f[45] >= `INH(p[98])) ? `INH(p[98]) : f[45];
        f[45] = (f[45] >= `INH(p[100])) ? `INH(p[100]) : f[45];
        f[45] = (f[45] > p[101]) ? p[101] : f[45];
        f[46] = 4095;
        f[46] = (f[46] > p[29]) ? p[29] : f[46];
        f[46] = (f[46] >= `INH(p[103])) ? `INH(p[103]) : f[46];
        f[47] = 4095;
        f[47] = (f[47] > p[102]) ? p[102] : f[47];
        f[47] = (f[47] >= `INH(p[104])) ? `INH(p[104]) : f[47];
        f[48] = 4095;
        f[48] = (f[48] >= `INH(p[29])) ? `INH(p[29]) : f[48];
        f[48] = (f[48] >= `INH(p[103])) ? `INH(p[103]) : f[48];
        f[48] = (f[48] > p[104]) ? p[104] : f[48];
        f[49] = 4095;
        f[49] = (f[49] >= `INH(p[102])) ? `INH(p[102]) : f[49];
        f[49] = (f[49] >= `INH(p[104])) ? `INH(p[104]) : f[49];
        f[49] = (f[49] > p[105]) ? p[105] : f[49];
        f[50] = 4095;
        f[50] = (f[50] >= `INH(p[0])) ? `INH(p[0]) : f[50];
        f[50] = (f[50] > p[99]) ? p[99] : f[50];
        f[50] = (f[50] > p[103]) ? p[103] : f[50];
        f[51] = 4095;
        f[51] = (f[51] > p[85]) ? p[85] : f[51];
        f[51] = (f[51] >= `INH(p[101])) ? `INH(p[101]) : f[51];
        f[51] = (f[51] >= `INH(p[105])) ? `INH(p[105]) : f[51];
        f[52] = 4095;
        f[52] = (f[52] > p[86]) ? p[86] : f[52];
        f[52] = (f[52] >= `INH(p[106])) ? `INH(p[106]) : f[52];
        f[53] = 4095;
        f[53] = (f[53] > p[30]) ? p[30] : f[53];
        f[53] = (f[53] >= `INH(p[87])) ? `INH(p[87]) : f[53];
        f[54] = 4095;
        f[54] = (f[54] >= `INH(p[30])) ? `INH(p[30]) : f[54];
        f[54] = (f[54] >= `INH(p[87])) ? `INH(p[87]) : f[54];
        f[54] = (f[54] > p[106]) ? p[106] : f[54];
        f[55] = 4095;
        f[55] = (f[55] > p[1]) ? p[1] : f[55];
        f[55] = (f[55] >= `INH(p[86])) ? `INH(p[86]) : f[55];
        f[55] = (f[55] >= `INH(p[106])) ? `INH(p[106]) : f[55];
        f[56] = 4095;
        f[56] = (f[56] >= `INH(p[108])) ? `INH(p[108]) : f[56];
        f[56] = (f[56] >= `INH(p[109])) ? `INH(p[109]) : f[56];
        f[56] = (f[56] > p[113]) ? p[113] : f[56];
        f[57] = 4095;
        f[57] = (f[57] > p[107]) ? p[107] : f[57];
        f[57] = (f[57] >= `INH(p[113])) ? `INH(p[113]) : f[57];
        f[58] = 4095;
        f[58] = (f[58] > p[111]) ? p[111] : f[58];
        f[58] = (f[58] >= `INH(p[113])) ? `INH(p[113]) : f[58];
        f[59] = 4095;
        f[59] = (f[59] >= p[108]/2) ? p[108]/2 : f[59];
        f[59] = (f[59] >= `INH(p[112])) ? `INH(p[112]) : f[59];
        f[60] = 4095;
        f[60] = (f[60] >= `INH(p[112])) ? `INH(p[112]) : f[60];
        f[60] = (f[60] > p[115]) ? p[115] : f[60];
        f[61] = 4095;
        f[61] = (f[61] > p[108]) ? p[108] : f[61];
        f[61] = (f[61] >= `INH(p[115])) ? `INH(p[115]) : f[61];
        f[61] = (f[61] > p[117]) ? p[117] : f[61];
        f[62] = 4095;
        f[62] = (f[62] >= `INH(p[115])) ? `INH(p[115]) : f[62];
        f[62] = (f[62] > p[118]) ? p[118] : f[62];
        f[63] = 4095;
        f[63] = (f[63] > p[107]) ? p[107] : f[63];
        f[63] = (f[63] >= `INH(p[117])) ? `INH(p[117]) : f[63];
        f[63] = (f[63] >= `INH(p[118])) ? `INH(p[118]) : f[63];
        f[64] = 4095;
        f[64] = (f[64] > p[107]) ? p[107] : f[64];
        f[64] = (f[64] >= `INH(p[116])) ? `INH(p[116]) : f[64];
        f[64] = (f[64] >= `INH(p[118])) ? `INH(p[118]) : f[64];
        f[65] = 4095;
        f[65] = (f[65] >= `INH(p[118])) ? `INH(p[118]) : f[65];
        f[65] = (f[65] > p[120]) ? p[120] : f[65];
        f[66] = 4095;
        f[66] = (f[66] > p[114]) ? p[114] : f[66];
        f[66] = (f[66] >= `INH(p[120])) ? `INH(p[120]) : f[66];
        f[67] = 4095;
        f[67] = (f[67] >= `INH(p[120])) ? `INH(p[120]) : f[67];
        f[67] = (f[67] > p[121]) ? p[121] : f[67];
        f[68] = 4095;
        f[68] = (f[68] > p[119]) ? p[119] : f[68];
        f[68] = (f[68] >= `INH(p[121])) ? `INH(p[121]) : f[68];
        f[69] = 4095;
        f[69] = (f[69] > p[109]) ? p[109] : f[69];
        f[69] = (f[69] > p[116]) ? p[116] : f[69];
        f[69] = (f[69] >= `INH(p[117])) ? `INH(p[117]) : f[69];
        f[69] = (f[69] >= `INH(p[121])) ? `INH(p[121]) : f[69];
        f[70] = 4095;
        f[70] = (f[70] > p[109]) ? p[109] : f[70];
        f[70] = (f[70] >= `INH(p[116])) ? `INH(p[116]) : f[70];
        f[70] = (f[70] >= `INH(p[121])) ? `INH(p[121]) : f[70];
        f[71] = 4095;
        f[71] = (f[71] > p[30]) ? p[30] : f[71];
        f[71] = (f[71] >= `INH(p[123])) ? `INH(p[123]) : f[71];
        f[72] = 4095;
        f[72] = (f[72] > p[122]) ? p[122] : f[72];
        f[72] = (f[72] >= `INH(p[124])) ? `INH(p[124]) : f[72];
        f[73] = 4095;
        f[73] = (f[73] >= `INH(p[30])) ? `INH(p[30]) : f[73];
        f[73] = (f[73] >= `INH(p[123])) ? `INH(p[123]) : f[73];
        f[73] = (f[73] > p[124]) ? p[124] : f[73];
        f[74] = 4095;
        f[74] = (f[74] >= `INH(p[122])) ? `INH(p[122]) : f[74];
        f[74] = (f[74] >= `INH(p[124])) ? `INH(p[124]) : f[74];
        f[74] = (f[74] > p[125]) ? p[125] : f[74];
        f[75] = 4095;
        f[75] = (f[75] > p[31]) ? p[31] : f[75];
        f[75] = (f[75] >= `INH(p[127])) ? `INH(p[127]) : f[75];
        f[76] = 4095;
        f[76] = (f[76] > p[126]) ? p[126] : f[76];
        f[76] = (f[76] >= `INH(p[128])) ? `INH(p[128]) : f[76];
        f[77] = 4095;
        f[77] = (f[77] >= `INH(p[31])) ? `INH(p[31]) : f[77];
        f[77] = (f[77] >= `INH(p[127])) ? `INH(p[127]) : f[77];
        f[77] = (f[77] > p[128]) ? p[128] : f[77];
        f[78] = 4095;
        f[78] = (f[78] >= `INH(p[126])) ? `INH(p[126]) : f[78];
        f[78] = (f[78] >= `INH(p[128])) ? `INH(p[128]) : f[78];
        f[78] = (f[78] > p[129]) ? p[129] : f[78];
        f[79] = 4095;
        f[79] = (f[79] >= `INH(p[1])) ? `INH(p[1]) : f[79];
        f[79] = (f[79] > p[123]) ? p[123] : f[79];
        f[79] = (f[79] > p[127]) ? p[127] : f[79];
        f[80] = 4095;
        f[80] = (f[80] > p[109]) ? p[109] : f[80];
        f[80] = (f[80] >= `INH(p[125])) ? `INH(p[125]) : f[80];
        f[80] = (f[80] >= `INH(p[129])) ? `INH(p[129]) : f[80];
        f[81] = 4095;
        f[81] = (f[81] > p[110]) ? p[110] : f[81];
        f[81] = (f[81] >= `INH(p[130])) ? `INH(p[130]) : f[81];
        f[82] = 4095;
        f[82] = (f[82] > p[32]) ? p[32] : f[82];
        f[82] = (f[82] >= `INH(p[111])) ? `INH(p[111]) : f[82];
        f[83] = 4095;
        f[83] = (f[83] >= `INH(p[32])) ? `INH(p[32]) : f[83];
        f[83] = (f[83] >= `INH(p[111])) ? `INH(p[111]) : f[83];
        f[83] = (f[83] > p[130]) ? p[130] : f[83];
        f[84] = 4095;
        f[84] = (f[84] > p[2]) ? p[2] : f[84];
        f[84] = (f[84] >= `INH(p[110])) ? `INH(p[110]) : f[84];
        f[84] = (f[84] >= `INH(p[130])) ? `INH(p[130]) : f[84];
        f[85] = 4095;
        f[85] = (f[85] >= `INH(p[132])) ? `INH(p[132]) : f[85];
        f[85] = (f[85] >= `INH(p[133])) ? `INH(p[133]) : f[85];
        f[85] = (f[85] > p[137]) ? p[137] : f[85];
        f[86] = 4095;
        f[86] = (f[86] > p[131]) ? p[131] : f[86];
        f[86] = (f[86] >= `INH(p[137])) ? `INH(p[137]) : f[86];
        f[87] = 4095;
        f[87] = (f[87] > p[135]) ? p[135] : f[87];
        f[87] = (f[87] >= `INH(p[137])) ? `INH(p[137]) : f[87];
        f[88] = 4095;
        f[88] = (f[88] >= p[132]/2) ? p[132]/2 : f[88];
        f[88] = (f[88] >= `INH(p[136])) ? `INH(p[136]) : f[88];
        f[89] = 4095;
        f[89] = (f[89] >= `INH(p[136])) ? `INH(p[136]) : f[89];
        f[89] = (f[89] > p[139]) ? p[139] : f[89];
        f[90] = 4095;
        f[90] = (f[90] > p[132]) ? p[132] : f[90];
        f[90] = (f[90] >= `INH(p[139])) ? `INH(p[139]) : f[90];
        f[90] = (f[90] > p[141]) ? p[141] : f[90];
        f[91] = 4095;
        f[91] = (f[91] >= `INH(p[139])) ? `INH(p[139]) : f[91];
        f[91] = (f[91] > p[142]) ? p[142] : f[91];
        f[92] = 4095;
        f[92] = (f[92] > p[131]) ? p[131] : f[92];
        f[92] = (f[92] >= `INH(p[141])) ? `INH(p[141]) : f[92];
        f[92] = (f[92] >= `INH(p[142])) ? `INH(p[142]) : f[92];
        f[93] = 4095;
        f[93] = (f[93] > p[131]) ? p[131] : f[93];
        f[93] = (f[93] >= `INH(p[140])) ? `INH(p[140]) : f[93];
        f[93] = (f[93] >= `INH(p[142])) ? `INH(p[142]) : f[93];
        f[94] = 4095;
        f[94] = (f[94] >= `INH(p[142])) ? `INH(p[142]) : f[94];
        f[94] = (f[94] > p[144]) ? p[144] : f[94];
        f[95] = 4095;
        f[95] = (f[95] > p[138]) ? p[138] : f[95];
        f[95] = (f[95] >= `INH(p[144])) ? `INH(p[144]) : f[95];
        f[96] = 4095;
        f[96] = (f[96] >= `INH(p[144])) ? `INH(p[144]) : f[96];
        f[96] = (f[96] > p[145]) ? p[145] : f[96];
        f[97] = 4095;
        f[97] = (f[97] > p[143]) ? p[143] : f[97];
        f[97] = (f[97] >= `INH(p[145])) ? `INH(p[145]) : f[97];
        f[98] = 4095;
        f[98] = (f[98] > p[133]) ? p[133] : f[98];
        f[98] = (f[98] > p[140]) ? p[140] : f[98];
        f[98] = (f[98] >= `INH(p[141])) ? `INH(p[141]) : f[98];
        f[98] = (f[98] >= `INH(p[145])) ? `INH(p[145]) : f[98];
        f[99] = 4095;
        f[99] = (f[99] > p[133]) ? p[133] : f[99];
        f[99] = (f[99] >= `INH(p[140])) ? `INH(p[140]) : f[99];
        f[99] = (f[99] >= `INH(p[145])) ? `INH(p[145]) : f[99];
        f[100] = 4095;
        f[100] = (f[100] > p[32]) ? p[32] : f[100];
        f[100] = (f[100] >= `INH(p[147])) ? `INH(p[147]) : f[100];
        f[101] = 4095;
        f[101] = (f[101] > p[146]) ? p[146] : f[101];
        f[101] = (f[101] >= `INH(p[148])) ? `INH(p[148]) : f[101];
        f[102] = 4095;
        f[102] = (f[102] >= `INH(p[32])) ? `INH(p[32]) : f[102];
        f[102] = (f[102] >= `INH(p[147])) ? `INH(p[147]) : f[102];
        f[102] = (f[102] > p[148]) ? p[148] : f[102];
        f[103] = 4095;
        f[103] = (f[103] >= `INH(p[146])) ? `INH(p[146]) : f[103];
        f[103] = (f[103] >= `INH(p[148])) ? `INH(p[148]) : f[103];
        f[103] = (f[103] > p[149]) ? p[149] : f[103];
        f[104] = 4095;
        f[104] = (f[104] > p[33]) ? p[33] : f[104];
        f[104] = (f[104] >= `INH(p[151])) ? `INH(p[151]) : f[104];
        f[105] = 4095;
        f[105] = (f[105] > p[150]) ? p[150] : f[105];
        f[105] = (f[105] >= `INH(p[152])) ? `INH(p[152]) : f[105];
        f[106] = 4095;
        f[106] = (f[106] >= `INH(p[33])) ? `INH(p[33]) : f[106];
        f[106] = (f[106] >= `INH(p[151])) ? `INH(p[151]) : f[106];
        f[106] = (f[106] > p[152]) ? p[152] : f[106];
        f[107] = 4095;
        f[107] = (f[107] >= `INH(p[150])) ? `INH(p[150]) : f[107];
        f[107] = (f[107] >= `INH(p[152])) ? `INH(p[152]) : f[107];
        f[107] = (f[107] > p[153]) ? p[153] : f[107];
        f[108] = 4095;
        f[108] = (f[108] >= `INH(p[2])) ? `INH(p[2]) : f[108];
        f[108] = (f[108] > p[147]) ? p[147] : f[108];
        f[108] = (f[108] > p[151]) ? p[151] : f[108];
        f[109] = 4095;
        f[109] = (f[109] > p[133]) ? p[133] : f[109];
        f[109] = (f[109] >= `INH(p[149])) ? `INH(p[149]) : f[109];
        f[109] = (f[109] >= `INH(p[153])) ? `INH(p[153]) : f[109];
        f[110] = 4095;
        f[110] = (f[110] > p[134]) ? p[134] : f[110];
        f[110] = (f[110] >= `INH(p[154])) ? `INH(p[154]) : f[110];
        f[111] = 4095;
        f[111] = (f[111] > p[34]) ? p[34] : f[111];
        f[111] = (f[111] >= `INH(p[135])) ? `INH(p[135]) : f[111];
        f[112] = 4095;
        f[112] = (f[112] >= `INH(p[34])) ? `INH(p[34]) : f[112];
        f[112] = (f[112] >= `INH(p[135])) ? `INH(p[135]) : f[112];
        f[112] = (f[112] > p[154]) ? p[154] : f[112];
        f[113] = 4095;
        f[113] = (f[113] > p[3]) ? p[3] : f[113];
        f[113] = (f[113] >= `INH(p[134])) ? `INH(p[134]) : f[113];
        f[113] = (f[113] >= `INH(p[154])) ? `INH(p[154]) : f[113];
        f[114] = 4095;
        f[114] = (f[114] >= `INH(p[156])) ? `INH(p[156]) : f[114];
        f[114] = (f[114] >= `INH(p[157])) ? `INH(p[157]) : f[114];
        f[114] = (f[114] > p[161]) ? p[161] : f[114];
        f[115] = 4095;
        f[115] = (f[115] > p[155]) ? p[155] : f[115];
        f[115] = (f[115] >= `INH(p[161])) ? `INH(p[161]) : f[115];
        f[116] = 4095;
        f[116] = (f[116] > p[159]) ? p[159] : f[116];
        f[116] = (f[116] >= `INH(p[161])) ? `INH(p[161]) : f[116];
        f[117] = 4095;
        f[117] = (f[117] >= p[156]/2) ? p[156]/2 : f[117];
        f[117] = (f[117] >= `INH(p[160])) ? `INH(p[160]) : f[117];
        f[118] = 4095;
        f[118] = (f[118] >= `INH(p[160])) ? `INH(p[160]) : f[118];
        f[118] = (f[118] > p[163]) ? p[163] : f[118];
        f[119] = 4095;
        f[119] = (f[119] > p[156]) ? p[156] : f[119];
        f[119] = (f[119] >= `INH(p[163])) ? `INH(p[163]) : f[119];
        f[119] = (f[119] > p[165]) ? p[165] : f[119];
        f[120] = 4095;
        f[120] = (f[120] >= `INH(p[163])) ? `INH(p[163]) : f[120];
        f[120] = (f[120] > p[166]) ? p[166] : f[120];
        f[121] = 4095;
        f[121] = (f[121] > p[155]) ? p[155] : f[121];
        f[121] = (f[121] >= `INH(p[165])) ? `INH(p[165]) : f[121];
        f[121] = (f[121] >= `INH(p[166])) ? `INH(p[166]) : f[121];
        f[122] = 4095;
        f[122] = (f[122] > p[155]) ? p[155] : f[122];
        f[122] = (f[122] >= `INH(p[164])) ? `INH(p[164]) : f[122];
        f[122] = (f[122] >= `INH(p[166])) ? `INH(p[166]) : f[122];
        f[123] = 4095;
        f[123] = (f[123] >= `INH(p[166])) ? `INH(p[166]) : f[123];
        f[123] = (f[123] > p[168]) ? p[168] : f[123];
        f[124] = 4095;
        f[124] = (f[124] > p[162]) ? p[162] : f[124];
        f[124] = (f[124] >= `INH(p[168])) ? `INH(p[168]) : f[124];
        f[125] = 4095;
        f[125] = (f[125] >= `INH(p[168])) ? `INH(p[168]) : f[125];
        f[125] = (f[125] > p[169]) ? p[169] : f[125];
        f[126] = 4095;
        f[126] = (f[126] > p[167]) ? p[167] : f[126];
        f[126] = (f[126] >= `INH(p[169])) ? `INH(p[169]) : f[126];
        f[127] = 4095;
        f[127] = (f[127] > p[157]) ? p[157] : f[127];
        f[127] = (f[127] > p[164]) ? p[164] : f[127];
        f[127] = (f[127] >= `INH(p[165])) ? `INH(p[165]) : f[127];
        f[127] = (f[127] >= `INH(p[169])) ? `INH(p[169]) : f[127];
        f[128] = 4095;
        f[128] = (f[128] > p[157]) ? p[157] : f[128];
        f[128] = (f[128] >= `INH(p[164])) ? `INH(p[164]) : f[128];
        f[128] = (f[128] >= `INH(p[169])) ? `INH(p[169]) : f[128];
        f[129] = 4095;
        f[129] = (f[129] > p[34]) ? p[34] : f[129];
        f[129] = (f[129] >= `INH(p[171])) ? `INH(p[171]) : f[129];
        f[130] = 4095;
        f[130] = (f[130] > p[170]) ? p[170] : f[130];
        f[130] = (f[130] >= `INH(p[172])) ? `INH(p[172]) : f[130];
        f[131] = 4095;
        f[131] = (f[131] >= `INH(p[34])) ? `INH(p[34]) : f[131];
        f[131] = (f[131] >= `INH(p[171])) ? `INH(p[171]) : f[131];
        f[131] = (f[131] > p[172]) ? p[172] : f[131];
        f[132] = 4095;
        f[132] = (f[132] >= `INH(p[170])) ? `INH(p[170]) : f[132];
        f[132] = (f[132] >= `INH(p[172])) ? `INH(p[172]) : f[132];
        f[132] = (f[132] > p[173]) ? p[173] : f[132];
        f[133] = 4095;
        f[133] = (f[133] > p[35]) ? p[35] : f[133];
        f[133] = (f[133] >= `INH(p[175])) ? `INH(p[175]) : f[133];
        f[134] = 4095;
        f[134] = (f[134] > p[174]) ? p[174] : f[134];
        f[134] = (f[134] >= `INH(p[176])) ? `INH(p[176]) : f[134];
        f[135] = 4095;
        f[135] = (f[135] >= `INH(p[35])) ? `INH(p[35]) : f[135];
        f[135] = (f[135] >= `INH(p[175])) ? `INH(p[175]) : f[135];
        f[135] = (f[135] > p[176]) ? p[176] : f[135];
        f[136] = 4095;
        f[136] = (f[136] >= `INH(p[174])) ? `INH(p[174]) : f[136];
        f[136] = (f[136] >= `INH(p[176])) ? `INH(p[176]) : f[136];
        f[136] = (f[136] > p[177]) ? p[177] : f[136];
        f[137] = 4095;
        f[137] = (f[137] >= `INH(p[3])) ? `INH(p[3]) : f[137];
        f[137] = (f[137] > p[171]) ? p[171] : f[137];
        f[137] = (f[137] > p[175]) ? p[175] : f[137];
        f[138] = 4095;
        f[138] = (f[138] > p[157]) ? p[157] : f[138];
        f[138] = (f[138] >= `INH(p[173])) ? `INH(p[173]) : f[138];
        f[138] = (f[138] >= `INH(p[177])) ? `INH(p[177]) : f[138];
        f[139] = 4095;
        f[139] = (f[139] > p[158]) ? p[158] : f[139];
        f[139] = (f[139] >= `INH(p[178])) ? `INH(p[178]) : f[139];
        f[140] = 4095;
        f[140] = (f[140] > p[36]) ? p[36] : f[140];
        f[140] = (f[140] >= `INH(p[159])) ? `INH(p[159]) : f[140];
        f[141] = 4095;
        f[141] = (f[141] >= `INH(p[36])) ? `INH(p[36]) : f[141];
        f[141] = (f[141] >= `INH(p[159])) ? `INH(p[159]) : f[141];
        f[141] = (f[141] > p[178]) ? p[178] : f[141];
        f[142] = 4095;
        f[142] = (f[142] > p[4]) ? p[4] : f[142];
        f[142] = (f[142] >= `INH(p[158])) ? `INH(p[158]) : f[142];
        f[142] = (f[142] >= `INH(p[178])) ? `INH(p[178]) : f[142];
        f[143] = 4095;
        f[143] = (f[143] >= `INH(p[180])) ? `INH(p[180]) : f[143];
        f[143] = (f[143] >= `INH(p[181])) ? `INH(p[181]) : f[143];
        f[143] = (f[143] > p[185]) ? p[185] : f[143];
        f[144] = 4095;
        f[144] = (f[144] > p[179]) ? p[179] : f[144];
        f[144] = (f[144] >= `INH(p[185])) ? `INH(p[185]) : f[144];
        f[145] = 4095;
        f[145] = (f[145] > p[183]) ? p[183] : f[145];
        f[145] = (f[145] >= `INH(p[185])) ? `INH(p[185]) : f[145];
        f[146] = 4095;
        f[146] = (f[146] >= p[180]/2) ? p[180]/2 : f[146];
        f[146] = (f[146] >= `INH(p[184])) ? `INH(p[184]) : f[146];
        f[147] = 4095;
        f[147] = (f[147] >= `INH(p[184])) ? `INH(p[184]) : f[147];
        f[147] = (f[147] > p[187]) ? p[187] : f[147];
        f[148] = 4095;
        f[148] = (f[148] > p[180]) ? p[180] : f[148];
        f[148] = (f[148] >= `INH(p[187])) ? `INH(p[187]) : f[148];
        f[148] = (f[148] > p[189]) ? p[189] : f[148];
        f[149] = 4095;
        f[149] = (f[149] >= `INH(p[187])) ? `INH(p[187]) : f[149];
        f[149] = (f[149] > p[190]) ? p[190] : f[149];
        f[150] = 4095;
        f[150] = (f[150] > p[179]) ? p[179] : f[150];
        f[150] = (f[150] >= `INH(p[189])) ? `INH(p[189]) : f[150];
        f[150] = (f[150] >= `INH(p[190])) ? `INH(p[190]) : f[150];
        f[151] = 4095;
        f[151] = (f[151] > p[179]) ? p[179] : f[151];
        f[151] = (f[151] >= `INH(p[188])) ? `INH(p[188]) : f[151];
        f[151] = (f[151] >= `INH(p[190])) ? `INH(p[190]) : f[151];
        f[152] = 4095;
        f[152] = (f[152] >= `INH(p[190])) ? `INH(p[190]) : f[152];
        f[152] = (f[152] > p[192]) ? p[192] : f[152];
        f[153] = 4095;
        f[153] = (f[153] > p[186]) ? p[186] : f[153];
        f[153] = (f[153] >= `INH(p[192])) ? `INH(p[192]) : f[153];
        f[154] = 4095;
        f[154] = (f[154] >= `INH(p[192])) ? `INH(p[192]) : f[154];
        f[154] = (f[154] > p[193]) ? p[193] : f[154];
        f[155] = 4095;
        f[155] = (f[155] > p[191]) ? p[191] : f[155];
        f[155] = (f[155] >= `INH(p[193])) ? `INH(p[193]) : f[155];
        f[156] = 4095;
        f[156] = (f[156] > p[181]) ? p[181] : f[156];
        f[156] = (f[156] > p[188]) ? p[188] : f[156];
        f[156] = (f[156] >= `INH(p[189])) ? `INH(p[189]) : f[156];
        f[156] = (f[156] >= `INH(p[193])) ? `INH(p[193]) : f[156];
        f[157] = 4095;
        f[157] = (f[157] > p[181]) ? p[181] : f[157];
        f[157] = (f[157] >= `INH(p[188])) ? `INH(p[188]) : f[157];
        f[157] = (f[157] >= `INH(p[193])) ? `INH(p[193]) : f[157];
        f[158] = 4095;
        f[158] = (f[158] > p[36]) ? p[36] : f[158];
        f[158] = (f[158] >= `INH(p[195])) ? `INH(p[195]) : f[158];
        f[159] = 4095;
        f[159] = (f[159] > p[194]) ? p[194] : f[159];
        f[159] = (f[159] >= `INH(p[196])) ? `INH(p[196]) : f[159];
        f[160] = 4095;
        f[160] = (f[160] >= `INH(p[36])) ? `INH(p[36]) : f[160];
        f[160] = (f[160] >= `INH(p[195])) ? `INH(p[195]) : f[160];
        f[160] = (f[160] > p[196]) ? p[196] : f[160];
        f[161] = 4095;
        f[161] = (f[161] >= `INH(p[194])) ? `INH(p[194]) : f[161];
        f[161] = (f[161] >= `INH(p[196])) ? `INH(p[196]) : f[161];
        f[161] = (f[161] > p[197]) ? p[197] : f[161];
        f[162] = 4095;
        f[162] = (f[162] > p[37]) ? p[37] : f[162];
        f[162] = (f[162] >= `INH(p[199])) ? `INH(p[199]) : f[162];
        f[163] = 4095;
        f[163] = (f[163] > p[198]) ? p[198] : f[163];
        f[163] = (f[163] >= `INH(p[200])) ? `INH(p[200]) : f[163];
        f[164] = 4095;
        f[164] = (f[164] >= `INH(p[37])) ? `INH(p[37]) : f[164];
        f[164] = (f[164] >= `INH(p[199])) ? `INH(p[199]) : f[164];
        f[164] = (f[164] > p[200]) ? p[200] : f[164];
        f[165] = 4095;
        f[165] = (f[165] >= `INH(p[198])) ? `INH(p[198]) : f[165];
        f[165] = (f[165] >= `INH(p[200])) ? `INH(p[200]) : f[165];
        f[165] = (f[165] > p[201]) ? p[201] : f[165];
        f[166] = 4095;
        f[166] = (f[166] >= `INH(p[4])) ? `INH(p[4]) : f[166];
        f[166] = (f[166] > p[195]) ? p[195] : f[166];
        f[166] = (f[166] > p[199]) ? p[199] : f[166];
        f[167] = 4095;
        f[167] = (f[167] > p[181]) ? p[181] : f[167];
        f[167] = (f[167] >= `INH(p[197])) ? `INH(p[197]) : f[167];
        f[167] = (f[167] >= `INH(p[201])) ? `INH(p[201]) : f[167];
        f[168] = 4095;
        f[168] = (f[168] > p[182]) ? p[182] : f[168];
        f[168] = (f[168] >= `INH(p[202])) ? `INH(p[202]) : f[168];
        f[169] = 4095;
        f[169] = (f[169] > p[38]) ? p[38] : f[169];
        f[169] = (f[169] >= `INH(p[183])) ? `INH(p[183]) : f[169];
        f[170] = 4095;
        f[170] = (f[170] >= `INH(p[38])) ? `INH(p[38]) : f[170];
        f[170] = (f[170] >= `INH(p[183])) ? `INH(p[183]) : f[170];
        f[170] = (f[170] > p[202]) ? p[202] : f[170];
        f[171] = 4095;
        f[171] = (f[171] > p[5]) ? p[5] : f[171];
        f[171] = (f[171] >= `INH(p[182])) ? `INH(p[182]) : f[171];
        f[171] = (f[171] >= `INH(p[202])) ? `INH(p[202]) : f[171];
        f[172] = 4095;
        f[172] = (f[172] >= `INH(p[204])) ? `INH(p[204]) : f[172];
        f[172] = (f[172] >= `INH(p[205])) ? `INH(p[205]) : f[172];
        f[172] = (f[172] > p[209]) ? p[209] : f[172];
        f[173] = 4095;
        f[173] = (f[173] > p[203]) ? p[203] : f[173];
        f[173] = (f[173] >= `INH(p[209])) ? `INH(p[209]) : f[173];
        f[174] = 4095;
        f[174] = (f[174] > p[207]) ? p[207] : f[174];
        f[174] = (f[174] >= `INH(p[209])) ? `INH(p[209]) : f[174];
        f[175] = 4095;
        f[175] = (f[175] >= p[204]/2) ? p[204]/2 : f[175];
        f[175] = (f[175] >= `INH(p[208])) ? `INH(p[208]) : f[175];
        f[176] = 4095;
        f[176] = (f[176] >= `INH(p[208])) ? `INH(p[208]) : f[176];
        f[176] = (f[176] > p[211]) ? p[211] : f[176];
        f[177] = 4095;
        f[177] = (f[177] > p[204]) ? p[204] : f[177];
        f[177] = (f[177] >= `INH(p[211])) ? `INH(p[211]) : f[177];
        f[177] = (f[177] > p[213]) ? p[213] : f[177];
        f[178] = 4095;
        f[178] = (f[178] >= `INH(p[211])) ? `INH(p[211]) : f[178];
        f[178] = (f[178] > p[214]) ? p[214] : f[178];
        f[179] = 4095;
        f[179] = (f[179] > p[203]) ? p[203] : f[179];
        f[179] = (f[179] >= `INH(p[213])) ? `INH(p[213]) : f[179];
        f[179] = (f[179] >= `INH(p[214])) ? `INH(p[214]) : f[179];
        f[180] = 4095;
        f[180] = (f[180] > p[203]) ? p[203] : f[180];
        f[180] = (f[180] >= `INH(p[212])) ? `INH(p[212]) : f[180];
        f[180] = (f[180] >= `INH(p[214])) ? `INH(p[214]) : f[180];
        f[181] = 4095;
        f[181] = (f[181] >= `INH(p[214])) ? `INH(p[214]) : f[181];
        f[181] = (f[181] > p[216]) ? p[216] : f[181];
        f[182] = 4095;
        f[182] = (f[182] > p[210]) ? p[210] : f[182];
        f[182] = (f[182] >= `INH(p[216])) ? `INH(p[216]) : f[182];
        f[183] = 4095;
        f[183] = (f[183] >= `INH(p[216])) ? `INH(p[216]) : f[183];
        f[183] = (f[183] > p[217]) ? p[217] : f[183];
        f[184] = 4095;
        f[184] = (f[184] > p[215]) ? p[215] : f[184];
        f[184] = (f[184] >= `INH(p[217])) ? `INH(p[217]) : f[184];
        f[185] = 4095;
        f[185] = (f[185] > p[205]) ? p[205] : f[185];
        f[185] = (f[185] > p[212]) ? p[212] : f[185];
        f[185] = (f[185] >= `INH(p[213])) ? `INH(p[213]) : f[185];
        f[185] = (f[185] >= `INH(p[217])) ? `INH(p[217]) : f[185];
        f[186] = 4095;
        f[186] = (f[186] > p[205]) ? p[205] : f[186];
        f[186] = (f[186] >= `INH(p[212])) ? `INH(p[212]) : f[186];
        f[186] = (f[186] >= `INH(p[217])) ? `INH(p[217]) : f[186];
        f[187] = 4095;
        f[187] = (f[187] > p[38]) ? p[38] : f[187];
        f[187] = (f[187] >= `INH(p[219])) ? `INH(p[219]) : f[187];
        f[188] = 4095;
        f[188] = (f[188] > p[218]) ? p[218] : f[188];
        f[188] = (f[188] >= `INH(p[220])) ? `INH(p[220]) : f[188];
        f[189] = 4095;
        f[189] = (f[189] >= `INH(p[38])) ? `INH(p[38]) : f[189];
        f[189] = (f[189] >= `INH(p[219])) ? `INH(p[219]) : f[189];
        f[189] = (f[189] > p[220]) ? p[220] : f[189];
        f[190] = 4095;
        f[190] = (f[190] >= `INH(p[218])) ? `INH(p[218]) : f[190];
        f[190] = (f[190] >= `INH(p[220])) ? `INH(p[220]) : f[190];
        f[190] = (f[190] > p[221]) ? p[221] : f[190];
        f[191] = 4095;
        f[191] = (f[191] > p[39]) ? p[39] : f[191];
        f[191] = (f[191] >= `INH(p[223])) ? `INH(p[223]) : f[191];
        f[192] = 4095;
        f[192] = (f[192] > p[222]) ? p[222] : f[192];
        f[192] = (f[192] >= `INH(p[224])) ? `INH(p[224]) : f[192];
        f[193] = 4095;
        f[193] = (f[193] >= `INH(p[39])) ? `INH(p[39]) : f[193];
        f[193] = (f[193] >= `INH(p[223])) ? `INH(p[223]) : f[193];
        f[193] = (f[193] > p[224]) ? p[224] : f[193];
        f[194] = 4095;
        f[194] = (f[194] >= `INH(p[222])) ? `INH(p[222]) : f[194];
        f[194] = (f[194] >= `INH(p[224])) ? `INH(p[224]) : f[194];
        f[194] = (f[194] > p[225]) ? p[225] : f[194];
        f[195] = 4095;
        f[195] = (f[195] >= `INH(p[5])) ? `INH(p[5]) : f[195];
        f[195] = (f[195] > p[219]) ? p[219] : f[195];
        f[195] = (f[195] > p[223]) ? p[223] : f[195];
        f[196] = 4095;
        f[196] = (f[196] > p[205]) ? p[205] : f[196];
        f[196] = (f[196] >= `INH(p[221])) ? `INH(p[221]) : f[196];
        f[196] = (f[196] >= `INH(p[225])) ? `INH(p[225]) : f[196];
        f[197] = 4095;
        f[197] = (f[197] > p[206]) ? p[206] : f[197];
        f[197] = (f[197] >= `INH(p[226])) ? `INH(p[226]) : f[197];
        f[198] = 4095;
        f[198] = (f[198] > p[40]) ? p[40] : f[198];
        f[198] = (f[198] >= `INH(p[207])) ? `INH(p[207]) : f[198];
        f[199] = 4095;
        f[199] = (f[199] >= `INH(p[40])) ? `INH(p[40]) : f[199];
        f[199] = (f[199] >= `INH(p[207])) ? `INH(p[207]) : f[199];
        f[199] = (f[199] > p[226]) ? p[226] : f[199];
        f[200] = 4095;
        f[200] = (f[200] > p[6]) ? p[6] : f[200];
        f[200] = (f[200] >= `INH(p[206])) ? `INH(p[206]) : f[200];
        f[200] = (f[200] >= `INH(p[226])) ? `INH(p[226]) : f[200];
        f[201] = 4095;
        f[201] = (f[201] >= `INH(p[228])) ? `INH(p[228]) : f[201];
        f[201] = (f[201] >= `INH(p[229])) ? `INH(p[229]) : f[201];
        f[201] = (f[201] > p[233]) ? p[233] : f[201];
        f[202] = 4095;
        f[202] = (f[202] > p[227]) ? p[227] : f[202];
        f[202] = (f[202] >= `INH(p[233])) ? `INH(p[233]) : f[202];
        f[203] = 4095;
        f[203] = (f[203] > p[231]) ? p[231] : f[203];
        f[203] = (f[203] >= `INH(p[233])) ? `INH(p[233]) : f[203];
        f[204] = 4095;
        f[204] = (f[204] >= p[228]/2) ? p[228]/2 : f[204];
        f[204] = (f[204] >= `INH(p[232])) ? `INH(p[232]) : f[204];
        f[205] = 4095;
        f[205] = (f[205] >= `INH(p[232])) ? `INH(p[232]) : f[205];
        f[205] = (f[205] > p[235]) ? p[235] : f[205];
        f[206] = 4095;
        f[206] = (f[206] > p[228]) ? p[228] : f[206];
        f[206] = (f[206] >= `INH(p[235])) ? `INH(p[235]) : f[206];
        f[206] = (f[206] > p[237]) ? p[237] : f[206];
        f[207] = 4095;
        f[207] = (f[207] >= `INH(p[235])) ? `INH(p[235]) : f[207];
        f[207] = (f[207] > p[238]) ? p[238] : f[207];
        f[208] = 4095;
        f[208] = (f[208] > p[227]) ? p[227] : f[208];
        f[208] = (f[208] >= `INH(p[237])) ? `INH(p[237]) : f[208];
        f[208] = (f[208] >= `INH(p[238])) ? `INH(p[238]) : f[208];
        f[209] = 4095;
        f[209] = (f[209] > p[227]) ? p[227] : f[209];
        f[209] = (f[209] >= `INH(p[236])) ? `INH(p[236]) : f[209];
        f[209] = (f[209] >= `INH(p[238])) ? `INH(p[238]) : f[209];
        f[210] = 4095;
        f[210] = (f[210] >= `INH(p[238])) ? `INH(p[238]) : f[210];
        f[210] = (f[210] > p[240]) ? p[240] : f[210];
        f[211] = 4095;
        f[211] = (f[211] > p[234]) ? p[234] : f[211];
        f[211] = (f[211] >= `INH(p[240])) ? `INH(p[240]) : f[211];
        f[212] = 4095;
        f[212] = (f[212] >= `INH(p[240])) ? `INH(p[240]) : f[212];
        f[212] = (f[212] > p[241]) ? p[241] : f[212];
        f[213] = 4095;
        f[213] = (f[213] > p[239]) ? p[239] : f[213];
        f[213] = (f[213] >= `INH(p[241])) ? `INH(p[241]) : f[213];
        f[214] = 4095;
        f[214] = (f[214] > p[229]) ? p[229] : f[214];
        f[214] = (f[214] > p[236]) ? p[236] : f[214];
        f[214] = (f[214] >= `INH(p[237])) ? `INH(p[237]) : f[214];
        f[214] = (f[214] >= `INH(p[241])) ? `INH(p[241]) : f[214];
        f[215] = 4095;
        f[215] = (f[215] > p[229]) ? p[229] : f[215];
        f[215] = (f[215] >= `INH(p[236])) ? `INH(p[236]) : f[215];
        f[215] = (f[215] >= `INH(p[241])) ? `INH(p[241]) : f[215];
        f[216] = 4095;
        f[216] = (f[216] > p[41]) ? p[41] : f[216];
        f[216] = (f[216] >= `INH(p[243])) ? `INH(p[243]) : f[216];
        f[217] = 4095;
        f[217] = (f[217] > p[242]) ? p[242] : f[217];
        f[217] = (f[217] >= `INH(p[244])) ? `INH(p[244]) : f[217];
        f[218] = 4095;
        f[218] = (f[218] >= `INH(p[41])) ? `INH(p[41]) : f[218];
        f[218] = (f[218] >= `INH(p[243])) ? `INH(p[243]) : f[218];
        f[218] = (f[218] > p[244]) ? p[244] : f[218];
        f[219] = 4095;
        f[219] = (f[219] >= `INH(p[242])) ? `INH(p[242]) : f[219];
        f[219] = (f[219] >= `INH(p[244])) ? `INH(p[244]) : f[219];
        f[219] = (f[219] > p[245]) ? p[245] : f[219];
        f[220] = 4095;
        f[220] = (f[220] > p[42]) ? p[42] : f[220];
        f[220] = (f[220] >= `INH(p[247])) ? `INH(p[247]) : f[220];
        f[221] = 4095;
        f[221] = (f[221] > p[246]) ? p[246] : f[221];
        f[221] = (f[221] >= `INH(p[248])) ? `INH(p[248]) : f[221];
        f[222] = 4095;
        f[222] = (f[222] >= `INH(p[42])) ? `INH(p[42]) : f[222];
        f[222] = (f[222] >= `INH(p[247])) ? `INH(p[247]) : f[222];
        f[222] = (f[222] > p[248]) ? p[248] : f[222];
        f[223] = 4095;
        f[223] = (f[223] >= `INH(p[246])) ? `INH(p[246]) : f[223];
        f[223] = (f[223] >= `INH(p[248])) ? `INH(p[248]) : f[223];
        f[223] = (f[223] > p[249]) ? p[249] : f[223];
        f[224] = 4095;
        f[224] = (f[224] >= `INH(p[6])) ? `INH(p[6]) : f[224];
        f[224] = (f[224] > p[243]) ? p[243] : f[224];
        f[224] = (f[224] > p[247]) ? p[247] : f[224];
        f[225] = 4095;
        f[225] = (f[225] > p[229]) ? p[229] : f[225];
        f[225] = (f[225] >= `INH(p[245])) ? `INH(p[245]) : f[225];
        f[225] = (f[225] >= `INH(p[249])) ? `INH(p[249]) : f[225];
        f[226] = 4095;
        f[226] = (f[226] > p[230]) ? p[230] : f[226];
        f[226] = (f[226] >= `INH(p[250])) ? `INH(p[250]) : f[226];
        f[227] = 4095;
        f[227] = (f[227] > p[43]) ? p[43] : f[227];
        f[227] = (f[227] >= `INH(p[231])) ? `INH(p[231]) : f[227];
        f[228] = 4095;
        f[228] = (f[228] >= `INH(p[43])) ? `INH(p[43]) : f[228];
        f[228] = (f[228] >= `INH(p[231])) ? `INH(p[231]) : f[228];
        f[228] = (f[228] > p[250]) ? p[250] : f[228];
        f[229] = 4095;
        f[229] = (f[229] > p[7]) ? p[7] : f[229];
        f[229] = (f[229] >= `INH(p[230])) ? `INH(p[230]) : f[229];
        f[229] = (f[229] >= `INH(p[250])) ? `INH(p[250]) : f[229];
        f[230] = 4095;
        f[230] = (f[230] >= `INH(p[252])) ? `INH(p[252]) : f[230];
        f[230] = (f[230] >= `INH(p[253])) ? `INH(p[253]) : f[230];
        f[230] = (f[230] > p[257]) ? p[257] : f[230];
        f[231] = 4095;
        f[231] = (f[231] > p[251]) ? p[251] : f[231];
        f[231] = (f[231] >= `INH(p[257])) ? `INH(p[257]) : f[231];
        f[232] = 4095;
        f[232] = (f[232] > p[255]) ? p[255] : f[232];
        f[232] = (f[232] >= `INH(p[257])) ? `INH(p[257]) : f[232];
        f[233] = 4095;
        f[233] = (f[233] >= p[252]/2) ? p[252]/2 : f[233];
        f[233] = (f[233] >= `INH(p[256])) ? `INH(p[256]) : f[233];
        f[234] = 4095;
        f[234] = (f[234] >= `INH(p[256])) ? `INH(p[256]) : f[234];
        f[234] = (f[234] > p[259]) ? p[259] : f[234];
        f[235] = 4095;
        f[235] = (f[235] > p[252]) ? p[252] : f[235];
        f[235] = (f[235] >= `INH(p[259])) ? `INH(p[259]) : f[235];
        f[235] = (f[235] > p[261]) ? p[261] : f[235];
        f[236] = 4095;
        f[236] = (f[236] >= `INH(p[259])) ? `INH(p[259]) : f[236];
        f[236] = (f[236] > p[262]) ? p[262] : f[236];
        f[237] = 4095;
        f[237] = (f[237] > p[251]) ? p[251] : f[237];
        f[237] = (f[237] >= `INH(p[261])) ? `INH(p[261]) : f[237];
        f[237] = (f[237] >= `INH(p[262])) ? `INH(p[262]) : f[237];
        f[238] = 4095;
        f[238] = (f[238] > p[251]) ? p[251] : f[238];
        f[238] = (f[238] >= `INH(p[260])) ? `INH(p[260]) : f[238];
        f[238] = (f[238] >= `INH(p[262])) ? `INH(p[262]) : f[238];
        f[239] = 4095;
        f[239] = (f[239] >= `INH(p[262])) ? `INH(p[262]) : f[239];
        f[239] = (f[239] > p[264]) ? p[264] : f[239];
        f[240] = 4095;
        f[240] = (f[240] > p[258]) ? p[258] : f[240];
        f[240] = (f[240] >= `INH(p[264])) ? `INH(p[264]) : f[240];
        f[241] = 4095;
        f[241] = (f[241] >= `INH(p[264])) ? `INH(p[264]) : f[241];
        f[241] = (f[241] > p[265]) ? p[265] : f[241];
        f[242] = 4095;
        f[242] = (f[242] > p[263]) ? p[263] : f[242];
        f[242] = (f[242] >= `INH(p[265])) ? `INH(p[265]) : f[242];
        f[243] = 4095;
        f[243] = (f[243] > p[253]) ? p[253] : f[243];
        f[243] = (f[243] > p[260]) ? p[260] : f[243];
        f[243] = (f[243] >= `INH(p[261])) ? `INH(p[261]) : f[243];
        f[243] = (f[243] >= `INH(p[265])) ? `INH(p[265]) : f[243];
        f[244] = 4095;
        f[244] = (f[244] > p[253]) ? p[253] : f[244];
        f[244] = (f[244] >= `INH(p[260])) ? `INH(p[260]) : f[244];
        f[244] = (f[244] >= `INH(p[265])) ? `INH(p[265]) : f[244];
        f[245] = 4095;
        f[245] = (f[245] > p[43]) ? p[43] : f[245];
        f[245] = (f[245] >= `INH(p[267])) ? `INH(p[267]) : f[245];
        f[246] = 4095;
        f[246] = (f[246] > p[266]) ? p[266] : f[246];
        f[246] = (f[246] >= `INH(p[268])) ? `INH(p[268]) : f[246];
        f[247] = 4095;
        f[247] = (f[247] >= `INH(p[43])) ? `INH(p[43]) : f[247];
        f[247] = (f[247] >= `INH(p[267])) ? `INH(p[267]) : f[247];
        f[247] = (f[247] > p[268]) ? p[268] : f[247];
        f[248] = 4095;
        f[248] = (f[248] >= `INH(p[266])) ? `INH(p[266]) : f[248];
        f[248] = (f[248] >= `INH(p[268])) ? `INH(p[268]) : f[248];
        f[248] = (f[248] > p[269]) ? p[269] : f[248];
        f[249] = 4095;
        f[249] = (f[249] > p[44]) ? p[44] : f[249];
        f[249] = (f[249] >= `INH(p[271])) ? `INH(p[271]) : f[249];
        f[250] = 4095;
        f[250] = (f[250] > p[270]) ? p[270] : f[250];
        f[250] = (f[250] >= `INH(p[272])) ? `INH(p[272]) : f[250];
        f[251] = 4095;
        f[251] = (f[251] >= `INH(p[44])) ? `INH(p[44]) : f[251];
        f[251] = (f[251] >= `INH(p[271])) ? `INH(p[271]) : f[251];
        f[251] = (f[251] > p[272]) ? p[272] : f[251];
        f[252] = 4095;
        f[252] = (f[252] >= `INH(p[270])) ? `INH(p[270]) : f[252];
        f[252] = (f[252] >= `INH(p[272])) ? `INH(p[272]) : f[252];
        f[252] = (f[252] > p[273]) ? p[273] : f[252];
        f[253] = 4095;
        f[253] = (f[253] >= `INH(p[7])) ? `INH(p[7]) : f[253];
        f[253] = (f[253] > p[267]) ? p[267] : f[253];
        f[253] = (f[253] > p[271]) ? p[271] : f[253];
        f[254] = 4095;
        f[254] = (f[254] > p[253]) ? p[253] : f[254];
        f[254] = (f[254] >= `INH(p[269])) ? `INH(p[269]) : f[254];
        f[254] = (f[254] >= `INH(p[273])) ? `INH(p[273]) : f[254];
        f[255] = 4095;
        f[255] = (f[255] > p[254]) ? p[254] : f[255];
        f[255] = (f[255] >= `INH(p[274])) ? `INH(p[274]) : f[255];
        f[256] = 4095;
        f[256] = (f[256] > p[45]) ? p[45] : f[256];
        f[256] = (f[256] >= `INH(p[255])) ? `INH(p[255]) : f[256];
        f[257] = 4095;
        f[257] = (f[257] >= `INH(p[45])) ? `INH(p[45]) : f[257];
        f[257] = (f[257] >= `INH(p[255])) ? `INH(p[255]) : f[257];
        f[257] = (f[257] > p[274]) ? p[274] : f[257];
        f[258] = 4095;
        f[258] = (f[258] > p[8]) ? p[8] : f[258];
        f[258] = (f[258] >= `INH(p[254])) ? `INH(p[254]) : f[258];
        f[258] = (f[258] >= `INH(p[274])) ? `INH(p[274]) : f[258];
        f[259] = 4095;
        f[259] = (f[259] >= `INH(p[276])) ? `INH(p[276]) : f[259];
        f[259] = (f[259] >= `INH(p[277])) ? `INH(p[277]) : f[259];
        f[259] = (f[259] > p[281]) ? p[281] : f[259];
        f[260] = 4095;
        f[260] = (f[260] > p[275]) ? p[275] : f[260];
        f[260] = (f[260] >= `INH(p[281])) ? `INH(p[281]) : f[260];
        f[261] = 4095;
        f[261] = (f[261] > p[279]) ? p[279] : f[261];
        f[261] = (f[261] >= `INH(p[281])) ? `INH(p[281]) : f[261];
        f[262] = 4095;
        f[262] = (f[262] >= p[276]/2) ? p[276]/2 : f[262];
        f[262] = (f[262] >= `INH(p[280])) ? `INH(p[280]) : f[262];
        f[263] = 4095;
        f[263] = (f[263] >= `INH(p[280])) ? `INH(p[280]) : f[263];
        f[263] = (f[263] > p[283]) ? p[283] : f[263];
        f[264] = 4095;
        f[264] = (f[264] > p[276]) ? p[276] : f[264];
        f[264] = (f[264] >= `INH(p[283])) ? `INH(p[283]) : f[264];
        f[264] = (f[264] > p[285]) ? p[285] : f[264];
        f[265] = 4095;
        f[265] = (f[265] >= `INH(p[283])) ? `INH(p[283]) : f[265];
        f[265] = (f[265] > p[286]) ? p[286] : f[265];
        f[266] = 4095;
        f[266] = (f[266] > p[275]) ? p[275] : f[266];
        f[266] = (f[266] >= `INH(p[285])) ? `INH(p[285]) : f[266];
        f[266] = (f[266] >= `INH(p[286])) ? `INH(p[286]) : f[266];
        f[267] = 4095;
        f[267] = (f[267] > p[275]) ? p[275] : f[267];
        f[267] = (f[267] >= `INH(p[284])) ? `INH(p[284]) : f[267];
        f[267] = (f[267] >= `INH(p[286])) ? `INH(p[286]) : f[267];
        f[268] = 4095;
        f[268] = (f[268] >= `INH(p[286])) ? `INH(p[286]) : f[268];
        f[268] = (f[268] > p[288]) ? p[288] : f[268];
        f[269] = 4095;
        f[269] = (f[269] > p[282]) ? p[282] : f[269];
        f[269] = (f[269] >= `INH(p[288])) ? `INH(p[288]) : f[269];
        f[270] = 4095;
        f[270] = (f[270] >= `INH(p[288])) ? `INH(p[288]) : f[270];
        f[270] = (f[270] > p[289]) ? p[289] : f[270];
        f[271] = 4095;
        f[271] = (f[271] > p[287]) ? p[287] : f[271];
        f[271] = (f[271] >= `INH(p[289])) ? `INH(p[289]) : f[271];
        f[272] = 4095;
        f[272] = (f[272] > p[277]) ? p[277] : f[272];
        f[272] = (f[272] > p[284]) ? p[284] : f[272];
        f[272] = (f[272] >= `INH(p[285])) ? `INH(p[285]) : f[272];
        f[272] = (f[272] >= `INH(p[289])) ? `INH(p[289]) : f[272];
        f[273] = 4095;
        f[273] = (f[273] > p[277]) ? p[277] : f[273];
        f[273] = (f[273] >= `INH(p[284])) ? `INH(p[284]) : f[273];
        f[273] = (f[273] >= `INH(p[289])) ? `INH(p[289]) : f[273];
        f[274] = 4095;
        f[274] = (f[274] > p[45]) ? p[45] : f[274];
        f[274] = (f[274] >= `INH(p[291])) ? `INH(p[291]) : f[274];
        f[275] = 4095;
        f[275] = (f[275] > p[290]) ? p[290] : f[275];
        f[275] = (f[275] >= `INH(p[292])) ? `INH(p[292]) : f[275];
        f[276] = 4095;
        f[276] = (f[276] >= `INH(p[45])) ? `INH(p[45]) : f[276];
        f[276] = (f[276] >= `INH(p[291])) ? `INH(p[291]) : f[276];
        f[276] = (f[276] > p[292]) ? p[292] : f[276];
        f[277] = 4095;
        f[277] = (f[277] >= `INH(p[290])) ? `INH(p[290]) : f[277];
        f[277] = (f[277] >= `INH(p[292])) ? `INH(p[292]) : f[277];
        f[277] = (f[277] > p[293]) ? p[293] : f[277];
        f[278] = 4095;
        f[278] = (f[278] > p[46]) ? p[46] : f[278];
        f[278] = (f[278] >= `INH(p[295])) ? `INH(p[295]) : f[278];
        f[279] = 4095;
        f[279] = (f[279] > p[294]) ? p[294] : f[279];
        f[279] = (f[279] >= `INH(p[296])) ? `INH(p[296]) : f[279];
        f[280] = 4095;
        f[280] = (f[280] >= `INH(p[46])) ? `INH(p[46]) : f[280];
        f[280] = (f[280] >= `INH(p[295])) ? `INH(p[295]) : f[280];
        f[280] = (f[280] > p[296]) ? p[296] : f[280];
        f[281] = 4095;
        f[281] = (f[281] >= `INH(p[294])) ? `INH(p[294]) : f[281];
        f[281] = (f[281] >= `INH(p[296])) ? `INH(p[296]) : f[281];
        f[281] = (f[281] > p[297]) ? p[297] : f[281];
        f[282] = 4095;
        f[282] = (f[282] >= `INH(p[8])) ? `INH(p[8]) : f[282];
        f[282] = (f[282] > p[291]) ? p[291] : f[282];
        f[282] = (f[282] > p[295]) ? p[295] : f[282];
        f[283] = 4095;
        f[283] = (f[283] > p[277]) ? p[277] : f[283];
        f[283] = (f[283] >= `INH(p[293])) ? `INH(p[293]) : f[283];
        f[283] = (f[283] >= `INH(p[297])) ? `INH(p[297]) : f[283];
        f[284] = 4095;
        f[284] = (f[284] > p[278]) ? p[278] : f[284];
        f[284] = (f[284] >= `INH(p[298])) ? `INH(p[298]) : f[284];
        f[285] = 4095;
        f[285] = (f[285] > p[47]) ? p[47] : f[285];
        f[285] = (f[285] >= `INH(p[279])) ? `INH(p[279]) : f[285];
        f[286] = 4095;
        f[286] = (f[286] >= `INH(p[47])) ? `INH(p[47]) : f[286];
        f[286] = (f[286] >= `INH(p[279])) ? `INH(p[279]) : f[286];
        f[286] = (f[286] > p[298]) ? p[298] : f[286];
        f[287] = 4095;
        f[287] = (f[287] > p[9]) ? p[9] : f[287];
        f[287] = (f[287] >= `INH(p[278])) ? `INH(p[278]) : f[287];
        f[287] = (f[287] >= `INH(p[298])) ? `INH(p[298]) : f[287];
        f[288] = 4095;
        f[288] = (f[288] >= `INH(p[300])) ? `INH(p[300]) : f[288];
        f[288] = (f[288] >= `INH(p[301])) ? `INH(p[301]) : f[288];
        f[288] = (f[288] > p[305]) ? p[305] : f[288];
        f[289] = 4095;
        f[289] = (f[289] > p[299]) ? p[299] : f[289];
        f[289] = (f[289] >= `INH(p[305])) ? `INH(p[305]) : f[289];
        f[290] = 4095;
        f[290] = (f[290] > p[303]) ? p[303] : f[290];
        f[290] = (f[290] >= `INH(p[305])) ? `INH(p[305]) : f[290];
        f[291] = 4095;
        f[291] = (f[291] >= p[300]/2) ? p[300]/2 : f[291];
        f[291] = (f[291] >= `INH(p[304])) ? `INH(p[304]) : f[291];
        f[292] = 4095;
        f[292] = (f[292] >= `INH(p[304])) ? `INH(p[304]) : f[292];
        f[292] = (f[292] > p[307]) ? p[307] : f[292];
        f[293] = 4095;
        f[293] = (f[293] > p[300]) ? p[300] : f[293];
        f[293] = (f[293] >= `INH(p[307])) ? `INH(p[307]) : f[293];
        f[293] = (f[293] > p[309]) ? p[309] : f[293];
        f[294] = 4095;
        f[294] = (f[294] >= `INH(p[307])) ? `INH(p[307]) : f[294];
        f[294] = (f[294] > p[310]) ? p[310] : f[294];
        f[295] = 4095;
        f[295] = (f[295] > p[299]) ? p[299] : f[295];
        f[295] = (f[295] >= `INH(p[309])) ? `INH(p[309]) : f[295];
        f[295] = (f[295] >= `INH(p[310])) ? `INH(p[310]) : f[295];
        f[296] = 4095;
        f[296] = (f[296] > p[299]) ? p[299] : f[296];
        f[296] = (f[296] >= `INH(p[308])) ? `INH(p[308]) : f[296];
        f[296] = (f[296] >= `INH(p[310])) ? `INH(p[310]) : f[296];
        f[297] = 4095;
        f[297] = (f[297] >= `INH(p[310])) ? `INH(p[310]) : f[297];
        f[297] = (f[297] > p[312]) ? p[312] : f[297];
        f[298] = 4095;
        f[298] = (f[298] > p[306]) ? p[306] : f[298];
        f[298] = (f[298] >= `INH(p[312])) ? `INH(p[312]) : f[298];
        f[299] = 4095;
        f[299] = (f[299] >= `INH(p[312])) ? `INH(p[312]) : f[299];
        f[299] = (f[299] > p[313]) ? p[313] : f[299];
        f[300] = 4095;
        f[300] = (f[300] > p[311]) ? p[311] : f[300];
        f[300] = (f[300] >= `INH(p[313])) ? `INH(p[313]) : f[300];
        f[301] = 4095;
        f[301] = (f[301] > p[301]) ? p[301] : f[301];
        f[301] = (f[301] > p[308]) ? p[308] : f[301];
        f[301] = (f[301] >= `INH(p[309])) ? `INH(p[309]) : f[301];
        f[301] = (f[301] >= `INH(p[313])) ? `INH(p[313]) : f[301];
        f[302] = 4095;
        f[302] = (f[302] > p[301]) ? p[301] : f[302];
        f[302] = (f[302] >= `INH(p[308])) ? `INH(p[308]) : f[302];
        f[302] = (f[302] >= `INH(p[313])) ? `INH(p[313]) : f[302];
        f[303] = 4095;
        f[303] = (f[303] > p[47]) ? p[47] : f[303];
        f[303] = (f[303] >= `INH(p[315])) ? `INH(p[315]) : f[303];
        f[304] = 4095;
        f[304] = (f[304] > p[314]) ? p[314] : f[304];
        f[304] = (f[304] >= `INH(p[316])) ? `INH(p[316]) : f[304];
        f[305] = 4095;
        f[305] = (f[305] >= `INH(p[47])) ? `INH(p[47]) : f[305];
        f[305] = (f[305] >= `INH(p[315])) ? `INH(p[315]) : f[305];
        f[305] = (f[305] > p[316]) ? p[316] : f[305];
        f[306] = 4095;
        f[306] = (f[306] >= `INH(p[314])) ? `INH(p[314]) : f[306];
        f[306] = (f[306] >= `INH(p[316])) ? `INH(p[316]) : f[306];
        f[306] = (f[306] > p[317]) ? p[317] : f[306];
        f[307] = 4095;
        f[307] = (f[307] > p[48]) ? p[48] : f[307];
        f[307] = (f[307] >= `INH(p[319])) ? `INH(p[319]) : f[307];
        f[308] = 4095;
        f[308] = (f[308] > p[318]) ? p[318] : f[308];
        f[308] = (f[308] >= `INH(p[320])) ? `INH(p[320]) : f[308];
        f[309] = 4095;
        f[309] = (f[309] >= `INH(p[48])) ? `INH(p[48]) : f[309];
        f[309] = (f[309] >= `INH(p[319])) ? `INH(p[319]) : f[309];
        f[309] = (f[309] > p[320]) ? p[320] : f[309];
        f[310] = 4095;
        f[310] = (f[310] >= `INH(p[318])) ? `INH(p[318]) : f[310];
        f[310] = (f[310] >= `INH(p[320])) ? `INH(p[320]) : f[310];
        f[310] = (f[310] > p[321]) ? p[321] : f[310];
        f[311] = 4095;
        f[311] = (f[311] >= `INH(p[9])) ? `INH(p[9]) : f[311];
        f[311] = (f[311] > p[315]) ? p[315] : f[311];
        f[311] = (f[311] > p[319]) ? p[319] : f[311];
        f[312] = 4095;
        f[312] = (f[312] > p[301]) ? p[301] : f[312];
        f[312] = (f[312] >= `INH(p[317])) ? `INH(p[317]) : f[312];
        f[312] = (f[312] >= `INH(p[321])) ? `INH(p[321]) : f[312];
        f[313] = 4095;
        f[313] = (f[313] > p[302]) ? p[302] : f[313];
        f[313] = (f[313] >= `INH(p[322])) ? `INH(p[322]) : f[313];
        f[314] = 4095;
        f[314] = (f[314] > p[49]) ? p[49] : f[314];
        f[314] = (f[314] >= `INH(p[303])) ? `INH(p[303]) : f[314];
        f[315] = 4095;
        f[315] = (f[315] >= `INH(p[49])) ? `INH(p[49]) : f[315];
        f[315] = (f[315] >= `INH(p[303])) ? `INH(p[303]) : f[315];
        f[315] = (f[315] > p[322]) ? p[322] : f[315];
        f[316] = 4095;
        f[316] = (f[316] > p[10]) ? p[10] : f[316];
        f[316] = (f[316] >= `INH(p[302])) ? `INH(p[302]) : f[316];
        f[316] = (f[316] >= `INH(p[322])) ? `INH(p[322]) : f[316];
        f[317] = 4095;
        f[317] = (f[317] >= `INH(p[324])) ? `INH(p[324]) : f[317];
        f[317] = (f[317] >= `INH(p[325])) ? `INH(p[325]) : f[317];
        f[317] = (f[317] > p[329]) ? p[329] : f[317];
        f[318] = 4095;
        f[318] = (f[318] > p[323]) ? p[323] : f[318];
        f[318] = (f[318] >= `INH(p[329])) ? `INH(p[329]) : f[318];
        f[319] = 4095;
        f[319] = (f[319] > p[327]) ? p[327] : f[319];
        f[319] = (f[319] >= `INH(p[329])) ? `INH(p[329]) : f[319];
        f[320] = 4095;
        f[320] = (f[320] >= p[324]/2) ? p[324]/2 : f[320];
        f[320] = (f[320] >= `INH(p[328])) ? `INH(p[328]) : f[320];
        f[321] = 4095;
        f[321] = (f[321] >= `INH(p[328])) ? `INH(p[328]) : f[321];
        f[321] = (f[321] > p[331]) ? p[331] : f[321];
        f[322] = 4095;
        f[322] = (f[322] > p[324]) ? p[324] : f[322];
        f[322] = (f[322] >= `INH(p[331])) ? `INH(p[331]) : f[322];
        f[322] = (f[322] > p[333]) ? p[333] : f[322];
        f[323] = 4095;
        f[323] = (f[323] >= `INH(p[331])) ? `INH(p[331]) : f[323];
        f[323] = (f[323] > p[334]) ? p[334] : f[323];
        f[324] = 4095;
        f[324] = (f[324] > p[323]) ? p[323] : f[324];
        f[324] = (f[324] >= `INH(p[333])) ? `INH(p[333]) : f[324];
        f[324] = (f[324] >= `INH(p[334])) ? `INH(p[334]) : f[324];
        f[325] = 4095;
        f[325] = (f[325] > p[323]) ? p[323] : f[325];
        f[325] = (f[325] >= `INH(p[332])) ? `INH(p[332]) : f[325];
        f[325] = (f[325] >= `INH(p[334])) ? `INH(p[334]) : f[325];
        f[326] = 4095;
        f[326] = (f[326] >= `INH(p[334])) ? `INH(p[334]) : f[326];
        f[326] = (f[326] > p[336]) ? p[336] : f[326];
        f[327] = 4095;
        f[327] = (f[327] > p[330]) ? p[330] : f[327];
        f[327] = (f[327] >= `INH(p[336])) ? `INH(p[336]) : f[327];
        f[328] = 4095;
        f[328] = (f[328] >= `INH(p[336])) ? `INH(p[336]) : f[328];
        f[328] = (f[328] > p[337]) ? p[337] : f[328];
        f[329] = 4095;
        f[329] = (f[329] > p[335]) ? p[335] : f[329];
        f[329] = (f[329] >= `INH(p[337])) ? `INH(p[337]) : f[329];
        f[330] = 4095;
        f[330] = (f[330] > p[325]) ? p[325] : f[330];
        f[330] = (f[330] > p[332]) ? p[332] : f[330];
        f[330] = (f[330] >= `INH(p[333])) ? `INH(p[333]) : f[330];
        f[330] = (f[330] >= `INH(p[337])) ? `INH(p[337]) : f[330];
        f[331] = 4095;
        f[331] = (f[331] > p[325]) ? p[325] : f[331];
        f[331] = (f[331] >= `INH(p[332])) ? `INH(p[332]) : f[331];
        f[331] = (f[331] >= `INH(p[337])) ? `INH(p[337]) : f[331];
        f[332] = 4095;
        f[332] = (f[332] > p[49]) ? p[49] : f[332];
        f[332] = (f[332] >= `INH(p[339])) ? `INH(p[339]) : f[332];
        f[333] = 4095;
        f[333] = (f[333] > p[338]) ? p[338] : f[333];
        f[333] = (f[333] >= `INH(p[340])) ? `INH(p[340]) : f[333];
        f[334] = 4095;
        f[334] = (f[334] >= `INH(p[49])) ? `INH(p[49]) : f[334];
        f[334] = (f[334] >= `INH(p[339])) ? `INH(p[339]) : f[334];
        f[334] = (f[334] > p[340]) ? p[340] : f[334];
        f[335] = 4095;
        f[335] = (f[335] >= `INH(p[338])) ? `INH(p[338]) : f[335];
        f[335] = (f[335] >= `INH(p[340])) ? `INH(p[340]) : f[335];
        f[335] = (f[335] > p[341]) ? p[341] : f[335];
        f[336] = 4095;
        f[336] = (f[336] > p[50]) ? p[50] : f[336];
        f[336] = (f[336] >= `INH(p[343])) ? `INH(p[343]) : f[336];
        f[337] = 4095;
        f[337] = (f[337] > p[342]) ? p[342] : f[337];
        f[337] = (f[337] >= `INH(p[344])) ? `INH(p[344]) : f[337];
        f[338] = 4095;
        f[338] = (f[338] >= `INH(p[50])) ? `INH(p[50]) : f[338];
        f[338] = (f[338] >= `INH(p[343])) ? `INH(p[343]) : f[338];
        f[338] = (f[338] > p[344]) ? p[344] : f[338];
        f[339] = 4095;
        f[339] = (f[339] >= `INH(p[342])) ? `INH(p[342]) : f[339];
        f[339] = (f[339] >= `INH(p[344])) ? `INH(p[344]) : f[339];
        f[339] = (f[339] > p[345]) ? p[345] : f[339];
        f[340] = 4095;
        f[340] = (f[340] >= `INH(p[10])) ? `INH(p[10]) : f[340];
        f[340] = (f[340] > p[339]) ? p[339] : f[340];
        f[340] = (f[340] > p[343]) ? p[343] : f[340];
        f[341] = 4095;
        f[341] = (f[341] > p[325]) ? p[325] : f[341];
        f[341] = (f[341] >= `INH(p[341])) ? `INH(p[341]) : f[341];
        f[341] = (f[341] >= `INH(p[345])) ? `INH(p[345]) : f[341];
        f[342] = 4095;
        f[342] = (f[342] > p[326]) ? p[326] : f[342];
        f[342] = (f[342] >= `INH(p[346])) ? `INH(p[346]) : f[342];
        f[343] = 4095;
        f[343] = (f[343] > p[51]) ? p[51] : f[343];
        f[343] = (f[343] >= `INH(p[327])) ? `INH(p[327]) : f[343];
        f[344] = 4095;
        f[344] = (f[344] >= `INH(p[51])) ? `INH(p[51]) : f[344];
        f[344] = (f[344] >= `INH(p[327])) ? `INH(p[327]) : f[344];
        f[344] = (f[344] > p[346]) ? p[346] : f[344];
        f[345] = 4095;
        f[345] = (f[345] > p[11]) ? p[11] : f[345];
        f[345] = (f[345] >= `INH(p[326])) ? `INH(p[326]) : f[345];
        f[345] = (f[345] >= `INH(p[346])) ? `INH(p[346]) : f[345];
        f[346] = 4095;
        f[346] = (f[346] > p[348]) ? p[348] : f[346];
        f[346] = (f[346] >= `INH(p[350])) ? `INH(p[350]) : f[346];
        f[347] = 4095;
        f[347] = (f[347] >= `INH(p[347])) ? `INH(p[347]) : f[347];
        f[347] = (f[347] >= `INH(p[348])) ? `INH(p[348]) : f[347];
        f[347] = (f[347] >= `INH(p[350])) ? `INH(p[350]) : f[347];
        f[347] = (f[347] > p[351]) ? p[351] : f[347];
        f[348] = 4095;
        f[348] = (f[348] > p[40]) ? p[40] : f[348];
        f[348] = (f[348] >= `INH(p[353])) ? `INH(p[353]) : f[348];
        f[349] = 4095;
        f[349] = (f[349] > p[352]) ? p[352] : f[349];
        f[349] = (f[349] >= `INH(p[354])) ? `INH(p[354]) : f[349];
        f[350] = 4095;
        f[350] = (f[350] >= `INH(p[40])) ? `INH(p[40]) : f[350];
        f[350] = (f[350] >= `INH(p[353])) ? `INH(p[353]) : f[350];
        f[350] = (f[350] > p[354]) ? p[354] : f[350];
        f[351] = 4095;
        f[351] = (f[351] >= `INH(p[352])) ? `INH(p[352]) : f[351];
        f[351] = (f[351] >= `INH(p[354])) ? `INH(p[354]) : f[351];
        f[351] = (f[351] > p[355]) ? p[355] : f[351];
        f[352] = 4095;
        f[352] = (f[352] > p[51]) ? p[51] : f[352];
        f[352] = (f[352] >= `INH(p[357])) ? `INH(p[357]) : f[352];
        f[353] = 4095;
        f[353] = (f[353] > p[356]) ? p[356] : f[353];
        f[353] = (f[353] >= `INH(p[358])) ? `INH(p[358]) : f[353];
        f[354] = 4095;
        f[354] = (f[354] >= `INH(p[51])) ? `INH(p[51]) : f[354];
        f[354] = (f[354] >= `INH(p[357])) ? `INH(p[357]) : f[354];
        f[354] = (f[354] > p[358]) ? p[358] : f[354];
        f[355] = 4095;
        f[355] = (f[355] >= `INH(p[356])) ? `INH(p[356]) : f[355];
        f[355] = (f[355] >= `INH(p[358])) ? `INH(p[358]) : f[355];
        f[355] = (f[355] > p[359]) ? p[359] : f[355];
        f[356] = 4095;
        f[356] = (f[356] >= `INH(p[11])) ? `INH(p[11]) : f[356];
        f[356] = (f[356] > p[353]) ? p[353] : f[356];
        f[356] = (f[356] > p[357]) ? p[357] : f[356];
        f[357] = 4095;
        f[357] = (f[357] > p[350]) ? p[350] : f[357];
        f[357] = (f[357] >= `INH(p[355])) ? `INH(p[355]) : f[357];
        f[357] = (f[357] >= `INH(p[359])) ? `INH(p[359]) : f[357];
        f[358] = 4095;
        f[358] = (f[358] > p[349]) ? p[349] : f[358];
        f[358] = (f[358] >= `INH(p[360])) ? `INH(p[360]) : f[358];
        f[359] = 4095;
        f[359] = (f[359] > p[52]) ? p[52] : f[359];
        f[359] = (f[359] >= `INH(p[351])) ? `INH(p[351]) : f[359];
        f[360] = 4095;
        f[360] = (f[360] >= `INH(p[52])) ? `INH(p[52]) : f[360];
        f[360] = (f[360] >= `INH(p[351])) ? `INH(p[351]) : f[360];
        f[360] = (f[360] > p[360]) ? p[360] : f[360];
        f[361] = 4095;
        f[361] = (f[361] > p[12]) ? p[12] : f[361];
        f[361] = (f[361] >= `INH(p[349])) ? `INH(p[349]) : f[361];
        f[361] = (f[361] >= `INH(p[360])) ? `INH(p[360]) : f[361];
        f[362] = 4095;
        f[362] = (f[362] >= `INH(p[362])) ? `INH(p[362]) : f[362];
        f[362] = (f[362] >= `INH(p[363])) ? `INH(p[363]) : f[362];
        f[362] = (f[362] > p[367]) ? p[367] : f[362];
        f[363] = 4095;
        f[363] = (f[363] > p[361]) ? p[361] : f[363];
        f[363] = (f[363] >= `INH(p[367])) ? `INH(p[367]) : f[363];
        f[364] = 4095;
        f[364] = (f[364] > p[365]) ? p[365] : f[364];
        f[364] = (f[364] >= `INH(p[367])) ? `INH(p[367]) : f[364];
        f[365] = 4095;
        f[365] = (f[365] >= p[362]/2) ? p[362]/2 : f[365];
        f[365] = (f[365] >= `INH(p[366])) ? `INH(p[366]) : f[365];
        f[366] = 4095;
        f[366] = (f[366] >= `INH(p[366])) ? `INH(p[366]) : f[366];
        f[366] = (f[366] > p[369]) ? p[369] : f[366];
        f[367] = 4095;
        f[367] = (f[367] > p[362]) ? p[362] : f[367];
        f[367] = (f[367] >= `INH(p[369])) ? `INH(p[369]) : f[367];
        f[367] = (f[367] > p[371]) ? p[371] : f[367];
        f[368] = 4095;
        f[368] = (f[368] >= `INH(p[369])) ? `INH(p[369]) : f[368];
        f[368] = (f[368] > p[372]) ? p[372] : f[368];
        f[369] = 4095;
        f[369] = (f[369] > p[361]) ? p[361] : f[369];
        f[369] = (f[369] >= `INH(p[371])) ? `INH(p[371]) : f[369];
        f[369] = (f[369] >= `INH(p[372])) ? `INH(p[372]) : f[369];
        f[370] = 4095;
        f[370] = (f[370] > p[361]) ? p[361] : f[370];
        f[370] = (f[370] >= `INH(p[370])) ? `INH(p[370]) : f[370];
        f[370] = (f[370] >= `INH(p[372])) ? `INH(p[372]) : f[370];
        f[371] = 4095;
        f[371] = (f[371] >= `INH(p[372])) ? `INH(p[372]) : f[371];
        f[371] = (f[371] > p[374]) ? p[374] : f[371];
        f[372] = 4095;
        f[372] = (f[372] > p[368]) ? p[368] : f[372];
        f[372] = (f[372] >= `INH(p[374])) ? `INH(p[374]) : f[372];
        f[373] = 4095;
        f[373] = (f[373] >= `INH(p[374])) ? `INH(p[374]) : f[373];
        f[373] = (f[373] > p[375]) ? p[375] : f[373];
        f[374] = 4095;
        f[374] = (f[374] > p[373]) ? p[373] : f[374];
        f[374] = (f[374] >= `INH(p[375])) ? `INH(p[375]) : f[374];
        f[375] = 4095;
        f[375] = (f[375] > p[363]) ? p[363] : f[375];
        f[375] = (f[375] > p[370]) ? p[370] : f[375];
        f[375] = (f[375] >= `INH(p[371])) ? `INH(p[371]) : f[375];
        f[375] = (f[375] >= `INH(p[375])) ? `INH(p[375]) : f[375];
        f[376] = 4095;
        f[376] = (f[376] > p[363]) ? p[363] : f[376];
        f[376] = (f[376] >= `INH(p[370])) ? `INH(p[370]) : f[376];
        f[376] = (f[376] >= `INH(p[375])) ? `INH(p[375]) : f[376];
        f[377] = 4095;
        f[377] = (f[377] > p[53]) ? p[53] : f[377];
        f[377] = (f[377] >= `INH(p[377])) ? `INH(p[377]) : f[377];
        f[378] = 4095;
        f[378] = (f[378] > p[376]) ? p[376] : f[378];
        f[378] = (f[378] >= `INH(p[378])) ? `INH(p[378]) : f[378];
        f[379] = 4095;
        f[379] = (f[379] >= `INH(p[53])) ? `INH(p[53]) : f[379];
        f[379] = (f[379] >= `INH(p[377])) ? `INH(p[377]) : f[379];
        f[379] = (f[379] > p[378]) ? p[378] : f[379];
        f[380] = 4095;
        f[380] = (f[380] >= `INH(p[376])) ? `INH(p[376]) : f[380];
        f[380] = (f[380] >= `INH(p[378])) ? `INH(p[378]) : f[380];
        f[380] = (f[380] > p[379]) ? p[379] : f[380];
        f[381] = 4095;
        f[381] = (f[381] > p[54]) ? p[54] : f[381];
        f[381] = (f[381] >= `INH(p[381])) ? `INH(p[381]) : f[381];
        f[382] = 4095;
        f[382] = (f[382] > p[380]) ? p[380] : f[382];
        f[382] = (f[382] >= `INH(p[382])) ? `INH(p[382]) : f[382];
        f[383] = 4095;
        f[383] = (f[383] >= `INH(p[54])) ? `INH(p[54]) : f[383];
        f[383] = (f[383] >= `INH(p[381])) ? `INH(p[381]) : f[383];
        f[383] = (f[383] > p[382]) ? p[382] : f[383];
        f[384] = 4095;
        f[384] = (f[384] >= `INH(p[380])) ? `INH(p[380]) : f[384];
        f[384] = (f[384] >= `INH(p[382])) ? `INH(p[382]) : f[384];
        f[384] = (f[384] > p[383]) ? p[383] : f[384];
        f[385] = 4095;
        f[385] = (f[385] >= `INH(p[12])) ? `INH(p[12]) : f[385];
        f[385] = (f[385] > p[377]) ? p[377] : f[385];
        f[385] = (f[385] > p[381]) ? p[381] : f[385];
        f[386] = 4095;
        f[386] = (f[386] > p[363]) ? p[363] : f[386];
        f[386] = (f[386] >= `INH(p[379])) ? `INH(p[379]) : f[386];
        f[386] = (f[386] >= `INH(p[383])) ? `INH(p[383]) : f[386];
        f[387] = 4095;
        f[387] = (f[387] > p[364]) ? p[364] : f[387];
        f[387] = (f[387] >= `INH(p[384])) ? `INH(p[384]) : f[387];
        f[388] = 4095;
        f[388] = (f[388] > p[55]) ? p[55] : f[388];
        f[388] = (f[388] >= `INH(p[365])) ? `INH(p[365]) : f[388];
        f[389] = 4095;
        f[389] = (f[389] >= `INH(p[55])) ? `INH(p[55]) : f[389];
        f[389] = (f[389] >= `INH(p[365])) ? `INH(p[365]) : f[389];
        f[389] = (f[389] > p[384]) ? p[384] : f[389];
        f[390] = 4095;
        f[390] = (f[390] > p[13]) ? p[13] : f[390];
        f[390] = (f[390] >= `INH(p[364])) ? `INH(p[364]) : f[390];
        f[390] = (f[390] >= `INH(p[384])) ? `INH(p[384]) : f[390];
        f[391] = 4095;
        f[391] = (f[391] >= `INH(p[386])) ? `INH(p[386]) : f[391];
        f[391] = (f[391] >= `INH(p[387])) ? `INH(p[387]) : f[391];
        f[391] = (f[391] > p[391]) ? p[391] : f[391];
        f[392] = 4095;
        f[392] = (f[392] > p[385]) ? p[385] : f[392];
        f[392] = (f[392] >= `INH(p[391])) ? `INH(p[391]) : f[392];
        f[393] = 4095;
        f[393] = (f[393] > p[389]) ? p[389] : f[393];
        f[393] = (f[393] >= `INH(p[391])) ? `INH(p[391]) : f[393];
        f[394] = 4095;
        f[394] = (f[394] >= p[386]/2) ? p[386]/2 : f[394];
        f[394] = (f[394] >= `INH(p[390])) ? `INH(p[390]) : f[394];
        f[395] = 4095;
        f[395] = (f[395] >= `INH(p[390])) ? `INH(p[390]) : f[395];
        f[395] = (f[395] > p[393]) ? p[393] : f[395];
        f[396] = 4095;
        f[396] = (f[396] > p[386]) ? p[386] : f[396];
        f[396] = (f[396] >= `INH(p[393])) ? `INH(p[393]) : f[396];
        f[396] = (f[396] > p[395]) ? p[395] : f[396];
        f[397] = 4095;
        f[397] = (f[397] >= `INH(p[393])) ? `INH(p[393]) : f[397];
        f[397] = (f[397] > p[396]) ? p[396] : f[397];
        f[398] = 4095;
        f[398] = (f[398] > p[385]) ? p[385] : f[398];
        f[398] = (f[398] >= `INH(p[395])) ? `INH(p[395]) : f[398];
        f[398] = (f[398] >= `INH(p[396])) ? `INH(p[396]) : f[398];
        f[399] = 4095;
        f[399] = (f[399] > p[385]) ? p[385] : f[399];
        f[399] = (f[399] >= `INH(p[394])) ? `INH(p[394]) : f[399];
        f[399] = (f[399] >= `INH(p[396])) ? `INH(p[396]) : f[399];
        f[400] = 4095;
        f[400] = (f[400] >= `INH(p[396])) ? `INH(p[396]) : f[400];
        f[400] = (f[400] > p[398]) ? p[398] : f[400];
        f[401] = 4095;
        f[401] = (f[401] > p[392]) ? p[392] : f[401];
        f[401] = (f[401] >= `INH(p[398])) ? `INH(p[398]) : f[401];
        f[402] = 4095;
        f[402] = (f[402] >= `INH(p[398])) ? `INH(p[398]) : f[402];
        f[402] = (f[402] > p[399]) ? p[399] : f[402];
        f[403] = 4095;
        f[403] = (f[403] > p[397]) ? p[397] : f[403];
        f[403] = (f[403] >= `INH(p[399])) ? `INH(p[399]) : f[403];
        f[404] = 4095;
        f[404] = (f[404] > p[387]) ? p[387] : f[404];
        f[404] = (f[404] > p[394]) ? p[394] : f[404];
        f[404] = (f[404] >= `INH(p[395])) ? `INH(p[395]) : f[404];
        f[404] = (f[404] >= `INH(p[399])) ? `INH(p[399]) : f[404];
        f[405] = 4095;
        f[405] = (f[405] > p[387]) ? p[387] : f[405];
        f[405] = (f[405] >= `INH(p[394])) ? `INH(p[394]) : f[405];
        f[405] = (f[405] >= `INH(p[399])) ? `INH(p[399]) : f[405];
        f[406] = 4095;
        f[406] = (f[406] > p[55]) ? p[55] : f[406];
        f[406] = (f[406] >= `INH(p[401])) ? `INH(p[401]) : f[406];
        f[407] = 4095;
        f[407] = (f[407] > p[400]) ? p[400] : f[407];
        f[407] = (f[407] >= `INH(p[402])) ? `INH(p[402]) : f[407];
        f[408] = 4095;
        f[408] = (f[408] >= `INH(p[55])) ? `INH(p[55]) : f[408];
        f[408] = (f[408] >= `INH(p[401])) ? `INH(p[401]) : f[408];
        f[408] = (f[408] > p[402]) ? p[402] : f[408];
        f[409] = 4095;
        f[409] = (f[409] >= `INH(p[400])) ? `INH(p[400]) : f[409];
        f[409] = (f[409] >= `INH(p[402])) ? `INH(p[402]) : f[409];
        f[409] = (f[409] > p[403]) ? p[403] : f[409];
        f[410] = 4095;
        f[410] = (f[410] > p[56]) ? p[56] : f[410];
        f[410] = (f[410] >= `INH(p[405])) ? `INH(p[405]) : f[410];
        f[411] = 4095;
        f[411] = (f[411] > p[404]) ? p[404] : f[411];
        f[411] = (f[411] >= `INH(p[406])) ? `INH(p[406]) : f[411];
        f[412] = 4095;
        f[412] = (f[412] >= `INH(p[56])) ? `INH(p[56]) : f[412];
        f[412] = (f[412] >= `INH(p[405])) ? `INH(p[405]) : f[412];
        f[412] = (f[412] > p[406]) ? p[406] : f[412];
        f[413] = 4095;
        f[413] = (f[413] >= `INH(p[404])) ? `INH(p[404]) : f[413];
        f[413] = (f[413] >= `INH(p[406])) ? `INH(p[406]) : f[413];
        f[413] = (f[413] > p[407]) ? p[407] : f[413];
        f[414] = 4095;
        f[414] = (f[414] >= `INH(p[13])) ? `INH(p[13]) : f[414];
        f[414] = (f[414] > p[401]) ? p[401] : f[414];
        f[414] = (f[414] > p[405]) ? p[405] : f[414];
        f[415] = 4095;
        f[415] = (f[415] > p[387]) ? p[387] : f[415];
        f[415] = (f[415] >= `INH(p[403])) ? `INH(p[403]) : f[415];
        f[415] = (f[415] >= `INH(p[407])) ? `INH(p[407]) : f[415];
        f[416] = 4095;
        f[416] = (f[416] > p[388]) ? p[388] : f[416];
        f[416] = (f[416] >= `INH(p[408])) ? `INH(p[408]) : f[416];
        f[417] = 4095;
        f[417] = (f[417] > p[57]) ? p[57] : f[417];
        f[417] = (f[417] >= `INH(p[389])) ? `INH(p[389]) : f[417];
        f[418] = 4095;
        f[418] = (f[418] >= `INH(p[57])) ? `INH(p[57]) : f[418];
        f[418] = (f[418] >= `INH(p[389])) ? `INH(p[389]) : f[418];
        f[418] = (f[418] > p[408]) ? p[408] : f[418];
        f[419] = 4095;
        f[419] = (f[419] > p[14]) ? p[14] : f[419];
        f[419] = (f[419] >= `INH(p[388])) ? `INH(p[388]) : f[419];
        f[419] = (f[419] >= `INH(p[408])) ? `INH(p[408]) : f[419];
        f[420] = 4095;
        f[420] = (f[420] >= `INH(p[410])) ? `INH(p[410]) : f[420];
        f[420] = (f[420] >= `INH(p[411])) ? `INH(p[411]) : f[420];
        f[420] = (f[420] > p[415]) ? p[415] : f[420];
        f[421] = 4095;
        f[421] = (f[421] > p[409]) ? p[409] : f[421];
        f[421] = (f[421] >= `INH(p[415])) ? `INH(p[415]) : f[421];
        f[422] = 4095;
        f[422] = (f[422] > p[413]) ? p[413] : f[422];
        f[422] = (f[422] >= `INH(p[415])) ? `INH(p[415]) : f[422];
        f[423] = 4095;
        f[423] = (f[423] >= p[410]/2) ? p[410]/2 : f[423];
        f[423] = (f[423] >= `INH(p[414])) ? `INH(p[414]) : f[423];
        f[424] = 4095;
        f[424] = (f[424] >= `INH(p[414])) ? `INH(p[414]) : f[424];
        f[424] = (f[424] > p[417]) ? p[417] : f[424];
        f[425] = 4095;
        f[425] = (f[425] > p[410]) ? p[410] : f[425];
        f[425] = (f[425] >= `INH(p[417])) ? `INH(p[417]) : f[425];
        f[425] = (f[425] > p[419]) ? p[419] : f[425];
        f[426] = 4095;
        f[426] = (f[426] >= `INH(p[417])) ? `INH(p[417]) : f[426];
        f[426] = (f[426] > p[420]) ? p[420] : f[426];
        f[427] = 4095;
        f[427] = (f[427] > p[409]) ? p[409] : f[427];
        f[427] = (f[427] >= `INH(p[419])) ? `INH(p[419]) : f[427];
        f[427] = (f[427] >= `INH(p[420])) ? `INH(p[420]) : f[427];
        f[428] = 4095;
        f[428] = (f[428] > p[409]) ? p[409] : f[428];
        f[428] = (f[428] >= `INH(p[418])) ? `INH(p[418]) : f[428];
        f[428] = (f[428] >= `INH(p[420])) ? `INH(p[420]) : f[428];
        f[429] = 4095;
        f[429] = (f[429] >= `INH(p[420])) ? `INH(p[420]) : f[429];
        f[429] = (f[429] > p[422]) ? p[422] : f[429];
        f[430] = 4095;
        f[430] = (f[430] > p[416]) ? p[416] : f[430];
        f[430] = (f[430] >= `INH(p[422])) ? `INH(p[422]) : f[430];
        f[431] = 4095;
        f[431] = (f[431] >= `INH(p[422])) ? `INH(p[422]) : f[431];
        f[431] = (f[431] > p[423]) ? p[423] : f[431];
        f[432] = 4095;
        f[432] = (f[432] > p[421]) ? p[421] : f[432];
        f[432] = (f[432] >= `INH(p[423])) ? `INH(p[423]) : f[432];
        f[433] = 4095;
        f[433] = (f[433] > p[411]) ? p[411] : f[433];
        f[433] = (f[433] > p[418]) ? p[418] : f[433];
        f[433] = (f[433] >= `INH(p[419])) ? `INH(p[419]) : f[433];
        f[433] = (f[433] >= `INH(p[423])) ? `INH(p[423]) : f[433];
        f[434] = 4095;
        f[434] = (f[434] > p[411]) ? p[411] : f[434];
        f[434] = (f[434] >= `INH(p[418])) ? `INH(p[418]) : f[434];
        f[434] = (f[434] >= `INH(p[423])) ? `INH(p[423]) : f[434];
        f[435] = 4095;
        f[435] = (f[435] > p[57]) ? p[57] : f[435];
        f[435] = (f[435] >= `INH(p[425])) ? `INH(p[425]) : f[435];
        f[436] = 4095;
        f[436] = (f[436] > p[424]) ? p[424] : f[436];
        f[436] = (f[436] >= `INH(p[426])) ? `INH(p[426]) : f[436];
        f[437] = 4095;
        f[437] = (f[437] >= `INH(p[57])) ? `INH(p[57]) : f[437];
        f[437] = (f[437] >= `INH(p[425])) ? `INH(p[425]) : f[437];
        f[437] = (f[437] > p[426]) ? p[426] : f[437];
        f[438] = 4095;
        f[438] = (f[438] >= `INH(p[424])) ? `INH(p[424]) : f[438];
        f[438] = (f[438] >= `INH(p[426])) ? `INH(p[426]) : f[438];
        f[438] = (f[438] > p[427]) ? p[427] : f[438];
        f[439] = 4095;
        f[439] = (f[439] > p[58]) ? p[58] : f[439];
        f[439] = (f[439] >= `INH(p[429])) ? `INH(p[429]) : f[439];
        f[440] = 4095;
        f[440] = (f[440] > p[428]) ? p[428] : f[440];
        f[440] = (f[440] >= `INH(p[430])) ? `INH(p[430]) : f[440];
        f[441] = 4095;
        f[441] = (f[441] >= `INH(p[58])) ? `INH(p[58]) : f[441];
        f[441] = (f[441] >= `INH(p[429])) ? `INH(p[429]) : f[441];
        f[441] = (f[441] > p[430]) ? p[430] : f[441];
        f[442] = 4095;
        f[442] = (f[442] >= `INH(p[428])) ? `INH(p[428]) : f[442];
        f[442] = (f[442] >= `INH(p[430])) ? `INH(p[430]) : f[442];
        f[442] = (f[442] > p[431]) ? p[431] : f[442];
        f[443] = 4095;
        f[443] = (f[443] >= `INH(p[14])) ? `INH(p[14]) : f[443];
        f[443] = (f[443] > p[425]) ? p[425] : f[443];
        f[443] = (f[443] > p[429]) ? p[429] : f[443];
        f[444] = 4095;
        f[444] = (f[444] > p[411]) ? p[411] : f[444];
        f[444] = (f[444] >= `INH(p[427])) ? `INH(p[427]) : f[444];
        f[444] = (f[444] >= `INH(p[431])) ? `INH(p[431]) : f[444];
        f[445] = 4095;
        f[445] = (f[445] > p[412]) ? p[412] : f[445];
        f[445] = (f[445] >= `INH(p[432])) ? `INH(p[432]) : f[445];
        f[446] = 4095;
        f[446] = (f[446] > p[59]) ? p[59] : f[446];
        f[446] = (f[446] >= `INH(p[413])) ? `INH(p[413]) : f[446];
        f[447] = 4095;
        f[447] = (f[447] >= `INH(p[59])) ? `INH(p[59]) : f[447];
        f[447] = (f[447] >= `INH(p[413])) ? `INH(p[413]) : f[447];
        f[447] = (f[447] > p[432]) ? p[432] : f[447];
        f[448] = 4095;
        f[448] = (f[448] > p[15]) ? p[15] : f[448];
        f[448] = (f[448] >= `INH(p[412])) ? `INH(p[412]) : f[448];
        f[448] = (f[448] >= `INH(p[432])) ? `INH(p[432]) : f[448];
        f[449] = 4095;
        f[449] = (f[449] >= `INH(p[434])) ? `INH(p[434]) : f[449];
        f[449] = (f[449] >= `INH(p[435])) ? `INH(p[435]) : f[449];
        f[449] = (f[449] > p[439]) ? p[439] : f[449];
        f[450] = 4095;
        f[450] = (f[450] > p[433]) ? p[433] : f[450];
        f[450] = (f[450] >= `INH(p[439])) ? `INH(p[439]) : f[450];
        f[451] = 4095;
        f[451] = (f[451] > p[437]) ? p[437] : f[451];
        f[451] = (f[451] >= `INH(p[439])) ? `INH(p[439]) : f[451];
        f[452] = 4095;
        f[452] = (f[452] >= p[434]/2) ? p[434]/2 : f[452];
        f[452] = (f[452] >= `INH(p[438])) ? `INH(p[438]) : f[452];
        f[453] = 4095;
        f[453] = (f[453] >= `INH(p[438])) ? `INH(p[438]) : f[453];
        f[453] = (f[453] > p[441]) ? p[441] : f[453];
        f[454] = 4095;
        f[454] = (f[454] > p[434]) ? p[434] : f[454];
        f[454] = (f[454] >= `INH(p[441])) ? `INH(p[441]) : f[454];
        f[454] = (f[454] > p[443]) ? p[443] : f[454];
        f[455] = 4095;
        f[455] = (f[455] >= `INH(p[441])) ? `INH(p[441]) : f[455];
        f[455] = (f[455] > p[444]) ? p[444] : f[455];
        f[456] = 4095;
        f[456] = (f[456] > p[433]) ? p[433] : f[456];
        f[456] = (f[456] >= `INH(p[443])) ? `INH(p[443]) : f[456];
        f[456] = (f[456] >= `INH(p[444])) ? `INH(p[444]) : f[456];
        f[457] = 4095;
        f[457] = (f[457] > p[433]) ? p[433] : f[457];
        f[457] = (f[457] >= `INH(p[442])) ? `INH(p[442]) : f[457];
        f[457] = (f[457] >= `INH(p[444])) ? `INH(p[444]) : f[457];
        f[458] = 4095;
        f[458] = (f[458] >= `INH(p[444])) ? `INH(p[444]) : f[458];
        f[458] = (f[458] > p[446]) ? p[446] : f[458];
        f[459] = 4095;
        f[459] = (f[459] > p[440]) ? p[440] : f[459];
        f[459] = (f[459] >= `INH(p[446])) ? `INH(p[446]) : f[459];
        f[460] = 4095;
        f[460] = (f[460] >= `INH(p[446])) ? `INH(p[446]) : f[460];
        f[460] = (f[460] > p[447]) ? p[447] : f[460];
        f[461] = 4095;
        f[461] = (f[461] > p[445]) ? p[445] : f[461];
        f[461] = (f[461] >= `INH(p[447])) ? `INH(p[447]) : f[461];
        f[462] = 4095;
        f[462] = (f[462] > p[435]) ? p[435] : f[462];
        f[462] = (f[462] > p[442]) ? p[442] : f[462];
        f[462] = (f[462] >= `INH(p[443])) ? `INH(p[443]) : f[462];
        f[462] = (f[462] >= `INH(p[447])) ? `INH(p[447]) : f[462];
        f[463] = 4095;
        f[463] = (f[463] > p[435]) ? p[435] : f[463];
        f[463] = (f[463] >= `INH(p[442])) ? `INH(p[442]) : f[463];
        f[463] = (f[463] >= `INH(p[447])) ? `INH(p[447]) : f[463];
        f[464] = 4095;
        f[464] = (f[464] > p[59]) ? p[59] : f[464];
        f[464] = (f[464] >= `INH(p[449])) ? `INH(p[449]) : f[464];
        f[465] = 4095;
        f[465] = (f[465] > p[448]) ? p[448] : f[465];
        f[465] = (f[465] >= `INH(p[450])) ? `INH(p[450]) : f[465];
        f[466] = 4095;
        f[466] = (f[466] >= `INH(p[59])) ? `INH(p[59]) : f[466];
        f[466] = (f[466] >= `INH(p[449])) ? `INH(p[449]) : f[466];
        f[466] = (f[466] > p[450]) ? p[450] : f[466];
        f[467] = 4095;
        f[467] = (f[467] >= `INH(p[448])) ? `INH(p[448]) : f[467];
        f[467] = (f[467] >= `INH(p[450])) ? `INH(p[450]) : f[467];
        f[467] = (f[467] > p[451]) ? p[451] : f[467];
        f[468] = 4095;
        f[468] = (f[468] > p[60]) ? p[60] : f[468];
        f[468] = (f[468] >= `INH(p[453])) ? `INH(p[453]) : f[468];
        f[469] = 4095;
        f[469] = (f[469] > p[452]) ? p[452] : f[469];
        f[469] = (f[469] >= `INH(p[454])) ? `INH(p[454]) : f[469];
        f[470] = 4095;
        f[470] = (f[470] >= `INH(p[60])) ? `INH(p[60]) : f[470];
        f[470] = (f[470] >= `INH(p[453])) ? `INH(p[453]) : f[470];
        f[470] = (f[470] > p[454]) ? p[454] : f[470];
        f[471] = 4095;
        f[471] = (f[471] >= `INH(p[452])) ? `INH(p[452]) : f[471];
        f[471] = (f[471] >= `INH(p[454])) ? `INH(p[454]) : f[471];
        f[471] = (f[471] > p[455]) ? p[455] : f[471];
        f[472] = 4095;
        f[472] = (f[472] >= `INH(p[15])) ? `INH(p[15]) : f[472];
        f[472] = (f[472] > p[449]) ? p[449] : f[472];
        f[472] = (f[472] > p[453]) ? p[453] : f[472];
        f[473] = 4095;
        f[473] = (f[473] > p[435]) ? p[435] : f[473];
        f[473] = (f[473] >= `INH(p[451])) ? `INH(p[451]) : f[473];
        f[473] = (f[473] >= `INH(p[455])) ? `INH(p[455]) : f[473];
        f[474] = 4095;
        f[474] = (f[474] > p[436]) ? p[436] : f[474];
        f[474] = (f[474] >= `INH(p[456])) ? `INH(p[456]) : f[474];
        f[475] = 4095;
        f[475] = (f[475] > p[61]) ? p[61] : f[475];
        f[475] = (f[475] >= `INH(p[437])) ? `INH(p[437]) : f[475];
        f[476] = 4095;
        f[476] = (f[476] >= `INH(p[61])) ? `INH(p[61]) : f[476];
        f[476] = (f[476] >= `INH(p[437])) ? `INH(p[437]) : f[476];
        f[476] = (f[476] > p[456]) ? p[456] : f[476];
        f[477] = 4095;
        f[477] = (f[477] > p[16]) ? p[16] : f[477];
        f[477] = (f[477] >= `INH(p[436])) ? `INH(p[436]) : f[477];
        f[477] = (f[477] >= `INH(p[456])) ? `INH(p[456]) : f[477];
        f[478] = 4095;
        f[478] = (f[478] > p[458]) ? p[458] : f[478];
        f[478] = (f[478] >= `INH(p[460])) ? `INH(p[460]) : f[478];
        f[479] = 4095;
        f[479] = (f[479] >= `INH(p[457])) ? `INH(p[457]) : f[479];
        f[479] = (f[479] >= `INH(p[458])) ? `INH(p[458]) : f[479];
        f[479] = (f[479] >= `INH(p[460])) ? `INH(p[460]) : f[479];
        f[479] = (f[479] > p[461]) ? p[461] : f[479];
        f[480] = 4095;
        f[480] = (f[480] > p[61]) ? p[61] : f[480];
        f[480] = (f[480] >= `INH(p[463])) ? `INH(p[463]) : f[480];
        f[481] = 4095;
        f[481] = (f[481] > p[462]) ? p[462] : f[481];
        f[481] = (f[481] >= `INH(p[464])) ? `INH(p[464]) : f[481];
        f[482] = 4095;
        f[482] = (f[482] >= `INH(p[61])) ? `INH(p[61]) : f[482];
        f[482] = (f[482] >= `INH(p[463])) ? `INH(p[463]) : f[482];
        f[482] = (f[482] > p[464]) ? p[464] : f[482];
        f[483] = 4095;
        f[483] = (f[483] >= `INH(p[462])) ? `INH(p[462]) : f[483];
        f[483] = (f[483] >= `INH(p[464])) ? `INH(p[464]) : f[483];
        f[483] = (f[483] > p[465]) ? p[465] : f[483];
        f[484] = 4095;
        f[484] = (f[484] > p[52]) ? p[52] : f[484];
        f[484] = (f[484] >= `INH(p[467])) ? `INH(p[467]) : f[484];
        f[485] = 4095;
        f[485] = (f[485] > p[466]) ? p[466] : f[485];
        f[485] = (f[485] >= `INH(p[468])) ? `INH(p[468]) : f[485];
        f[486] = 4095;
        f[486] = (f[486] >= `INH(p[52])) ? `INH(p[52]) : f[486];
        f[486] = (f[486] >= `INH(p[467])) ? `INH(p[467]) : f[486];
        f[486] = (f[486] > p[468]) ? p[468] : f[486];
        f[487] = 4095;
        f[487] = (f[487] >= `INH(p[466])) ? `INH(p[466]) : f[487];
        f[487] = (f[487] >= `INH(p[468])) ? `INH(p[468]) : f[487];
        f[487] = (f[487] > p[469]) ? p[469] : f[487];
        f[488] = 4095;
        f[488] = (f[488] >= `INH(p[16])) ? `INH(p[16]) : f[488];
        f[488] = (f[488] > p[463]) ? p[463] : f[488];
        f[488] = (f[488] > p[467]) ? p[467] : f[488];
        f[489] = 4095;
        f[489] = (f[489] > p[460]) ? p[460] : f[489];
        f[489] = (f[489] >= `INH(p[465])) ? `INH(p[465]) : f[489];
        f[489] = (f[489] >= `INH(p[469])) ? `INH(p[469]) : f[489];
        f[490] = 4095;
        f[490] = (f[490] > p[459]) ? p[459] : f[490];
        f[490] = (f[490] >= `INH(p[470])) ? `INH(p[470]) : f[490];
        f[491] = 4095;
        f[491] = (f[491] > p[62]) ? p[62] : f[491];
        f[491] = (f[491] >= `INH(p[461])) ? `INH(p[461]) : f[491];
        f[492] = 4095;
        f[492] = (f[492] >= `INH(p[62])) ? `INH(p[62]) : f[492];
        f[492] = (f[492] >= `INH(p[461])) ? `INH(p[461]) : f[492];
        f[492] = (f[492] > p[470]) ? p[470] : f[492];
        f[493] = 4095;
        f[493] = (f[493] > p[17]) ? p[17] : f[493];
        f[493] = (f[493] >= `INH(p[459])) ? `INH(p[459]) : f[493];
        f[493] = (f[493] >= `INH(p[470])) ? `INH(p[470]) : f[493];
        f[494] = 4095;
        f[494] = (f[494] >= `INH(p[472])) ? `INH(p[472]) : f[494];
        f[494] = (f[494] >= `INH(p[473])) ? `INH(p[473]) : f[494];
        f[494] = (f[494] > p[477]) ? p[477] : f[494];
        f[495] = 4095;
        f[495] = (f[495] > p[471]) ? p[471] : f[495];
        f[495] = (f[495] >= `INH(p[477])) ? `INH(p[477]) : f[495];
        f[496] = 4095;
        f[496] = (f[496] > p[475]) ? p[475] : f[496];
        f[496] = (f[496] >= `INH(p[477])) ? `INH(p[477]) : f[496];
        f[497] = 4095;
        f[497] = (f[497] >= p[472]/2) ? p[472]/2 : f[497];
        f[497] = (f[497] >= `INH(p[476])) ? `INH(p[476]) : f[497];
        f[498] = 4095;
        f[498] = (f[498] >= `INH(p[476])) ? `INH(p[476]) : f[498];
        f[498] = (f[498] > p[479]) ? p[479] : f[498];
        f[499] = 4095;
        f[499] = (f[499] > p[472]) ? p[472] : f[499];
        f[499] = (f[499] >= `INH(p[479])) ? `INH(p[479]) : f[499];
        f[499] = (f[499] > p[481]) ? p[481] : f[499];
        f[500] = 4095;
        f[500] = (f[500] >= `INH(p[479])) ? `INH(p[479]) : f[500];
        f[500] = (f[500] > p[482]) ? p[482] : f[500];
        f[501] = 4095;
        f[501] = (f[501] > p[471]) ? p[471] : f[501];
        f[501] = (f[501] >= `INH(p[481])) ? `INH(p[481]) : f[501];
        f[501] = (f[501] >= `INH(p[482])) ? `INH(p[482]) : f[501];
        f[502] = 4095;
        f[502] = (f[502] > p[471]) ? p[471] : f[502];
        f[502] = (f[502] >= `INH(p[480])) ? `INH(p[480]) : f[502];
        f[502] = (f[502] >= `INH(p[482])) ? `INH(p[482]) : f[502];
        f[503] = 4095;
        f[503] = (f[503] >= `INH(p[482])) ? `INH(p[482]) : f[503];
        f[503] = (f[503] > p[484]) ? p[484] : f[503];
        f[504] = 4095;
        f[504] = (f[504] > p[478]) ? p[478] : f[504];
        f[504] = (f[504] >= `INH(p[484])) ? `INH(p[484]) : f[504];
        f[505] = 4095;
        f[505] = (f[505] >= `INH(p[484])) ? `INH(p[484]) : f[505];
        f[505] = (f[505] > p[485]) ? p[485] : f[505];
        f[506] = 4095;
        f[506] = (f[506] > p[483]) ? p[483] : f[506];
        f[506] = (f[506] >= `INH(p[485])) ? `INH(p[485]) : f[506];
        f[507] = 4095;
        f[507] = (f[507] > p[473]) ? p[473] : f[507];
        f[507] = (f[507] > p[480]) ? p[480] : f[507];
        f[507] = (f[507] >= `INH(p[481])) ? `INH(p[481]) : f[507];
        f[507] = (f[507] >= `INH(p[485])) ? `INH(p[485]) : f[507];
        f[508] = 4095;
        f[508] = (f[508] > p[473]) ? p[473] : f[508];
        f[508] = (f[508] >= `INH(p[480])) ? `INH(p[480]) : f[508];
        f[508] = (f[508] >= `INH(p[485])) ? `INH(p[485]) : f[508];
        f[509] = 4095;
        f[509] = (f[509] > p[63]) ? p[63] : f[509];
        f[509] = (f[509] >= `INH(p[487])) ? `INH(p[487]) : f[509];
        f[510] = 4095;
        f[510] = (f[510] > p[486]) ? p[486] : f[510];
        f[510] = (f[510] >= `INH(p[488])) ? `INH(p[488]) : f[510];
        f[511] = 4095;
        f[511] = (f[511] >= `INH(p[63])) ? `INH(p[63]) : f[511];
        f[511] = (f[511] >= `INH(p[487])) ? `INH(p[487]) : f[511];
        f[511] = (f[511] > p[488]) ? p[488] : f[511];
        f[512] = 4095;
        f[512] = (f[512] >= `INH(p[486])) ? `INH(p[486]) : f[512];
        f[512] = (f[512] >= `INH(p[488])) ? `INH(p[488]) : f[512];
        f[512] = (f[512] > p[489]) ? p[489] : f[512];
        f[513] = 4095;
        f[513] = (f[513] > p[64]) ? p[64] : f[513];
        f[513] = (f[513] >= `INH(p[491])) ? `INH(p[491]) : f[513];
        f[514] = 4095;
        f[514] = (f[514] > p[490]) ? p[490] : f[514];
        f[514] = (f[514] >= `INH(p[492])) ? `INH(p[492]) : f[514];
        f[515] = 4095;
        f[515] = (f[515] >= `INH(p[64])) ? `INH(p[64]) : f[515];
        f[515] = (f[515] >= `INH(p[491])) ? `INH(p[491]) : f[515];
        f[515] = (f[515] > p[492]) ? p[492] : f[515];
        f[516] = 4095;
        f[516] = (f[516] >= `INH(p[490])) ? `INH(p[490]) : f[516];
        f[516] = (f[516] >= `INH(p[492])) ? `INH(p[492]) : f[516];
        f[516] = (f[516] > p[493]) ? p[493] : f[516];
        f[517] = 4095;
        f[517] = (f[517] >= `INH(p[17])) ? `INH(p[17]) : f[517];
        f[517] = (f[517] > p[487]) ? p[487] : f[517];
        f[517] = (f[517] > p[491]) ? p[491] : f[517];
        f[518] = 4095;
        f[518] = (f[518] > p[473]) ? p[473] : f[518];
        f[518] = (f[518] >= `INH(p[489])) ? `INH(p[489]) : f[518];
        f[518] = (f[518] >= `INH(p[493])) ? `INH(p[493]) : f[518];
        f[519] = 4095;
        f[519] = (f[519] > p[474]) ? p[474] : f[519];
        f[519] = (f[519] >= `INH(p[494])) ? `INH(p[494]) : f[519];
        f[520] = 4095;
        f[520] = (f[520] > p[65]) ? p[65] : f[520];
        f[520] = (f[520] >= `INH(p[475])) ? `INH(p[475]) : f[520];
        f[521] = 4095;
        f[521] = (f[521] >= `INH(p[65])) ? `INH(p[65]) : f[521];
        f[521] = (f[521] >= `INH(p[475])) ? `INH(p[475]) : f[521];
        f[521] = (f[521] > p[494]) ? p[494] : f[521];
        f[522] = 4095;
        f[522] = (f[522] > p[18]) ? p[18] : f[522];
        f[522] = (f[522] >= `INH(p[474])) ? `INH(p[474]) : f[522];
        f[522] = (f[522] >= `INH(p[494])) ? `INH(p[494]) : f[522];
        f[523] = 4095;
        f[523] = (f[523] >= `INH(p[496])) ? `INH(p[496]) : f[523];
        f[523] = (f[523] >= `INH(p[497])) ? `INH(p[497]) : f[523];
        f[523] = (f[523] > p[501]) ? p[501] : f[523];
        f[524] = 4095;
        f[524] = (f[524] > p[495]) ? p[495] : f[524];
        f[524] = (f[524] >= `INH(p[501])) ? `INH(p[501]) : f[524];
        f[525] = 4095;
        f[525] = (f[525] > p[499]) ? p[499] : f[525];
        f[525] = (f[525] >= `INH(p[501])) ? `INH(p[501]) : f[525];
        f[526] = 4095;
        f[526] = (f[526] >= p[496]/2) ? p[496]/2 : f[526];
        f[526] = (f[526] >= `INH(p[500])) ? `INH(p[500]) : f[526];
        f[527] = 4095;
        f[527] = (f[527] >= `INH(p[500])) ? `INH(p[500]) : f[527];
        f[527] = (f[527] > p[503]) ? p[503] : f[527];
        f[528] = 4095;
        f[528] = (f[528] > p[496]) ? p[496] : f[528];
        f[528] = (f[528] >= `INH(p[503])) ? `INH(p[503]) : f[528];
        f[528] = (f[528] > p[505]) ? p[505] : f[528];
        f[529] = 4095;
        f[529] = (f[529] >= `INH(p[503])) ? `INH(p[503]) : f[529];
        f[529] = (f[529] > p[506]) ? p[506] : f[529];
        f[530] = 4095;
        f[530] = (f[530] > p[495]) ? p[495] : f[530];
        f[530] = (f[530] >= `INH(p[505])) ? `INH(p[505]) : f[530];
        f[530] = (f[530] >= `INH(p[506])) ? `INH(p[506]) : f[530];
        f[531] = 4095;
        f[531] = (f[531] > p[495]) ? p[495] : f[531];
        f[531] = (f[531] >= `INH(p[504])) ? `INH(p[504]) : f[531];
        f[531] = (f[531] >= `INH(p[506])) ? `INH(p[506]) : f[531];
        f[532] = 4095;
        f[532] = (f[532] >= `INH(p[506])) ? `INH(p[506]) : f[532];
        f[532] = (f[532] > p[508]) ? p[508] : f[532];
        f[533] = 4095;
        f[533] = (f[533] > p[502]) ? p[502] : f[533];
        f[533] = (f[533] >= `INH(p[508])) ? `INH(p[508]) : f[533];
        f[534] = 4095;
        f[534] = (f[534] >= `INH(p[508])) ? `INH(p[508]) : f[534];
        f[534] = (f[534] > p[509]) ? p[509] : f[534];
        f[535] = 4095;
        f[535] = (f[535] > p[507]) ? p[507] : f[535];
        f[535] = (f[535] >= `INH(p[509])) ? `INH(p[509]) : f[535];
        f[536] = 4095;
        f[536] = (f[536] > p[497]) ? p[497] : f[536];
        f[536] = (f[536] > p[504]) ? p[504] : f[536];
        f[536] = (f[536] >= `INH(p[505])) ? `INH(p[505]) : f[536];
        f[536] = (f[536] >= `INH(p[509])) ? `INH(p[509]) : f[536];
        f[537] = 4095;
        f[537] = (f[537] > p[497]) ? p[497] : f[537];
        f[537] = (f[537] >= `INH(p[504])) ? `INH(p[504]) : f[537];
        f[537] = (f[537] >= `INH(p[509])) ? `INH(p[509]) : f[537];
        f[538] = 4095;
        f[538] = (f[538] > p[65]) ? p[65] : f[538];
        f[538] = (f[538] >= `INH(p[511])) ? `INH(p[511]) : f[538];
        f[539] = 4095;
        f[539] = (f[539] > p[510]) ? p[510] : f[539];
        f[539] = (f[539] >= `INH(p[512])) ? `INH(p[512]) : f[539];
        f[540] = 4095;
        f[540] = (f[540] >= `INH(p[65])) ? `INH(p[65]) : f[540];
        f[540] = (f[540] >= `INH(p[511])) ? `INH(p[511]) : f[540];
        f[540] = (f[540] > p[512]) ? p[512] : f[540];
        f[541] = 4095;
        f[541] = (f[541] >= `INH(p[510])) ? `INH(p[510]) : f[541];
        f[541] = (f[541] >= `INH(p[512])) ? `INH(p[512]) : f[541];
        f[541] = (f[541] > p[513]) ? p[513] : f[541];
        f[542] = 4095;
        f[542] = (f[542] > p[66]) ? p[66] : f[542];
        f[542] = (f[542] >= `INH(p[515])) ? `INH(p[515]) : f[542];
        f[543] = 4095;
        f[543] = (f[543] > p[514]) ? p[514] : f[543];
        f[543] = (f[543] >= `INH(p[516])) ? `INH(p[516]) : f[543];
        f[544] = 4095;
        f[544] = (f[544] >= `INH(p[66])) ? `INH(p[66]) : f[544];
        f[544] = (f[544] >= `INH(p[515])) ? `INH(p[515]) : f[544];
        f[544] = (f[544] > p[516]) ? p[516] : f[544];
        f[545] = 4095;
        f[545] = (f[545] >= `INH(p[514])) ? `INH(p[514]) : f[545];
        f[545] = (f[545] >= `INH(p[516])) ? `INH(p[516]) : f[545];
        f[545] = (f[545] > p[517]) ? p[517] : f[545];
        f[546] = 4095;
        f[546] = (f[546] >= `INH(p[18])) ? `INH(p[18]) : f[546];
        f[546] = (f[546] > p[511]) ? p[511] : f[546];
        f[546] = (f[546] > p[515]) ? p[515] : f[546];
        f[547] = 4095;
        f[547] = (f[547] > p[497]) ? p[497] : f[547];
        f[547] = (f[547] >= `INH(p[513])) ? `INH(p[513]) : f[547];
        f[547] = (f[547] >= `INH(p[517])) ? `INH(p[517]) : f[547];
        f[548] = 4095;
        f[548] = (f[548] > p[498]) ? p[498] : f[548];
        f[548] = (f[548] >= `INH(p[518])) ? `INH(p[518]) : f[548];
        f[549] = 4095;
        f[549] = (f[549] > p[67]) ? p[67] : f[549];
        f[549] = (f[549] >= `INH(p[499])) ? `INH(p[499]) : f[549];
        f[550] = 4095;
        f[550] = (f[550] >= `INH(p[67])) ? `INH(p[67]) : f[550];
        f[550] = (f[550] >= `INH(p[499])) ? `INH(p[499]) : f[550];
        f[550] = (f[550] > p[518]) ? p[518] : f[550];
        f[551] = 4095;
        f[551] = (f[551] > p[19]) ? p[19] : f[551];
        f[551] = (f[551] >= `INH(p[498])) ? `INH(p[498]) : f[551];
        f[551] = (f[551] >= `INH(p[518])) ? `INH(p[518]) : f[551];
        f[552] = 4095;
        f[552] = (f[552] >= `INH(p[520])) ? `INH(p[520]) : f[552];
        f[552] = (f[552] >= `INH(p[521])) ? `INH(p[521]) : f[552];
        f[552] = (f[552] > p[525]) ? p[525] : f[552];
        f[553] = 4095;
        f[553] = (f[553] > p[519]) ? p[519] : f[553];
        f[553] = (f[553] >= `INH(p[525])) ? `INH(p[525]) : f[553];
        f[554] = 4095;
        f[554] = (f[554] > p[523]) ? p[523] : f[554];
        f[554] = (f[554] >= `INH(p[525])) ? `INH(p[525]) : f[554];
        f[555] = 4095;
        f[555] = (f[555] >= p[520]/2) ? p[520]/2 : f[555];
        f[555] = (f[555] >= `INH(p[524])) ? `INH(p[524]) : f[555];
        f[556] = 4095;
        f[556] = (f[556] >= `INH(p[524])) ? `INH(p[524]) : f[556];
        f[556] = (f[556] > p[527]) ? p[527] : f[556];
        f[557] = 4095;
        f[557] = (f[557] > p[520]) ? p[520] : f[557];
        f[557] = (f[557] >= `INH(p[527])) ? `INH(p[527]) : f[557];
        f[557] = (f[557] > p[529]) ? p[529] : f[557];
        f[558] = 4095;
        f[558] = (f[558] >= `INH(p[527])) ? `INH(p[527]) : f[558];
        f[558] = (f[558] > p[530]) ? p[530] : f[558];
        f[559] = 4095;
        f[559] = (f[559] > p[519]) ? p[519] : f[559];
        f[559] = (f[559] >= `INH(p[529])) ? `INH(p[529]) : f[559];
        f[559] = (f[559] >= `INH(p[530])) ? `INH(p[530]) : f[559];
        f[560] = 4095;
        f[560] = (f[560] > p[519]) ? p[519] : f[560];
        f[560] = (f[560] >= `INH(p[528])) ? `INH(p[528]) : f[560];
        f[560] = (f[560] >= `INH(p[530])) ? `INH(p[530]) : f[560];
        f[561] = 4095;
        f[561] = (f[561] >= `INH(p[530])) ? `INH(p[530]) : f[561];
        f[561] = (f[561] > p[532]) ? p[532] : f[561];
        f[562] = 4095;
        f[562] = (f[562] > p[526]) ? p[526] : f[562];
        f[562] = (f[562] >= `INH(p[532])) ? `INH(p[532]) : f[562];
        f[563] = 4095;
        f[563] = (f[563] >= `INH(p[532])) ? `INH(p[532]) : f[563];
        f[563] = (f[563] > p[533]) ? p[533] : f[563];
        f[564] = 4095;
        f[564] = (f[564] > p[531]) ? p[531] : f[564];
        f[564] = (f[564] >= `INH(p[533])) ? `INH(p[533]) : f[564];
        f[565] = 4095;
        f[565] = (f[565] > p[521]) ? p[521] : f[565];
        f[565] = (f[565] > p[528]) ? p[528] : f[565];
        f[565] = (f[565] >= `INH(p[529])) ? `INH(p[529]) : f[565];
        f[565] = (f[565] >= `INH(p[533])) ? `INH(p[533]) : f[565];
        f[566] = 4095;
        f[566] = (f[566] > p[521]) ? p[521] : f[566];
        f[566] = (f[566] >= `INH(p[528])) ? `INH(p[528]) : f[566];
        f[566] = (f[566] >= `INH(p[533])) ? `INH(p[533]) : f[566];
        f[567] = 4095;
        f[567] = (f[567] > p[67]) ? p[67] : f[567];
        f[567] = (f[567] >= `INH(p[535])) ? `INH(p[535]) : f[567];
        f[568] = 4095;
        f[568] = (f[568] > p[534]) ? p[534] : f[568];
        f[568] = (f[568] >= `INH(p[536])) ? `INH(p[536]) : f[568];
        f[569] = 4095;
        f[569] = (f[569] >= `INH(p[67])) ? `INH(p[67]) : f[569];
        f[569] = (f[569] >= `INH(p[535])) ? `INH(p[535]) : f[569];
        f[569] = (f[569] > p[536]) ? p[536] : f[569];
        f[570] = 4095;
        f[570] = (f[570] >= `INH(p[534])) ? `INH(p[534]) : f[570];
        f[570] = (f[570] >= `INH(p[536])) ? `INH(p[536]) : f[570];
        f[570] = (f[570] > p[537]) ? p[537] : f[570];
        f[571] = 4095;
        f[571] = (f[571] > p[68]) ? p[68] : f[571];
        f[571] = (f[571] >= `INH(p[539])) ? `INH(p[539]) : f[571];
        f[572] = 4095;
        f[572] = (f[572] > p[538]) ? p[538] : f[572];
        f[572] = (f[572] >= `INH(p[540])) ? `INH(p[540]) : f[572];
        f[573] = 4095;
        f[573] = (f[573] >= `INH(p[68])) ? `INH(p[68]) : f[573];
        f[573] = (f[573] >= `INH(p[539])) ? `INH(p[539]) : f[573];
        f[573] = (f[573] > p[540]) ? p[540] : f[573];
        f[574] = 4095;
        f[574] = (f[574] >= `INH(p[538])) ? `INH(p[538]) : f[574];
        f[574] = (f[574] >= `INH(p[540])) ? `INH(p[540]) : f[574];
        f[574] = (f[574] > p[541]) ? p[541] : f[574];
        f[575] = 4095;
        f[575] = (f[575] >= `INH(p[19])) ? `INH(p[19]) : f[575];
        f[575] = (f[575] > p[535]) ? p[535] : f[575];
        f[575] = (f[575] > p[539]) ? p[539] : f[575];
        f[576] = 4095;
        f[576] = (f[576] > p[521]) ? p[521] : f[576];
        f[576] = (f[576] >= `INH(p[537])) ? `INH(p[537]) : f[576];
        f[576] = (f[576] >= `INH(p[541])) ? `INH(p[541]) : f[576];
        f[577] = 4095;
        f[577] = (f[577] > p[522]) ? p[522] : f[577];
        f[577] = (f[577] >= `INH(p[542])) ? `INH(p[542]) : f[577];
        f[578] = 4095;
        f[578] = (f[578] > p[69]) ? p[69] : f[578];
        f[578] = (f[578] >= `INH(p[523])) ? `INH(p[523]) : f[578];
        f[579] = 4095;
        f[579] = (f[579] >= `INH(p[69])) ? `INH(p[69]) : f[579];
        f[579] = (f[579] >= `INH(p[523])) ? `INH(p[523]) : f[579];
        f[579] = (f[579] > p[542]) ? p[542] : f[579];
        f[580] = 4095;
        f[580] = (f[580] > p[20]) ? p[20] : f[580];
        f[580] = (f[580] >= `INH(p[522])) ? `INH(p[522]) : f[580];
        f[580] = (f[580] >= `INH(p[542])) ? `INH(p[542]) : f[580];
        f[581] = 4095;
        f[581] = (f[581] > p[544]) ? p[544] : f[581];
        f[581] = (f[581] >= `INH(p[546])) ? `INH(p[546]) : f[581];
        f[582] = 4095;
        f[582] = (f[582] >= `INH(p[543])) ? `INH(p[543]) : f[582];
        f[582] = (f[582] >= `INH(p[544])) ? `INH(p[544]) : f[582];
        f[582] = (f[582] >= `INH(p[546])) ? `INH(p[546]) : f[582];
        f[582] = (f[582] > p[547]) ? p[547] : f[582];
        f[583] = 4095;
        f[583] = (f[583] > p[69]) ? p[69] : f[583];
        f[583] = (f[583] >= `INH(p[549])) ? `INH(p[549]) : f[583];
        f[584] = 4095;
        f[584] = (f[584] > p[548]) ? p[548] : f[584];
        f[584] = (f[584] >= `INH(p[550])) ? `INH(p[550]) : f[584];
        f[585] = 4095;
        f[585] = (f[585] >= `INH(p[69])) ? `INH(p[69]) : f[585];
        f[585] = (f[585] >= `INH(p[549])) ? `INH(p[549]) : f[585];
        f[585] = (f[585] > p[550]) ? p[550] : f[585];
        f[586] = 4095;
        f[586] = (f[586] >= `INH(p[548])) ? `INH(p[548]) : f[586];
        f[586] = (f[586] >= `INH(p[550])) ? `INH(p[550]) : f[586];
        f[586] = (f[586] > p[551]) ? p[551] : f[586];
        f[587] = 4095;
        f[587] = (f[587] > p[62]) ? p[62] : f[587];
        f[587] = (f[587] >= `INH(p[553])) ? `INH(p[553]) : f[587];
        f[588] = 4095;
        f[588] = (f[588] > p[552]) ? p[552] : f[588];
        f[588] = (f[588] >= `INH(p[554])) ? `INH(p[554]) : f[588];
        f[589] = 4095;
        f[589] = (f[589] >= `INH(p[62])) ? `INH(p[62]) : f[589];
        f[589] = (f[589] >= `INH(p[553])) ? `INH(p[553]) : f[589];
        f[589] = (f[589] > p[554]) ? p[554] : f[589];
        f[590] = 4095;
        f[590] = (f[590] >= `INH(p[552])) ? `INH(p[552]) : f[590];
        f[590] = (f[590] >= `INH(p[554])) ? `INH(p[554]) : f[590];
        f[590] = (f[590] > p[555]) ? p[555] : f[590];
        f[591] = 4095;
        f[591] = (f[591] >= `INH(p[20])) ? `INH(p[20]) : f[591];
        f[591] = (f[591] > p[549]) ? p[549] : f[591];
        f[591] = (f[591] > p[553]) ? p[553] : f[591];
        f[592] = 4095;
        f[592] = (f[592] > p[546]) ? p[546] : f[592];
        f[592] = (f[592] >= `INH(p[551])) ? `INH(p[551]) : f[592];
        f[592] = (f[592] >= `INH(p[555])) ? `INH(p[555]) : f[592];
        f[593] = 4095;
        f[593] = (f[593] > p[545]) ? p[545] : f[593];
        f[593] = (f[593] >= `INH(p[556])) ? `INH(p[556]) : f[593];
        f[594] = 4095;
        f[594] = (f[594] > p[70]) ? p[70] : f[594];
        f[594] = (f[594] >= `INH(p[547])) ? `INH(p[547]) : f[594];
        f[595] = 4095;
        f[595] = (f[595] >= `INH(p[70])) ? `INH(p[70]) : f[595];
        f[595] = (f[595] >= `INH(p[547])) ? `INH(p[547]) : f[595];
        f[595] = (f[595] > p[556]) ? p[556] : f[595];
        f[596] = 4095;
        f[596] = (f[596] > p[21]) ? p[21] : f[596];
        f[596] = (f[596] >= `INH(p[545])) ? `INH(p[545]) : f[596];
        f[596] = (f[596] >= `INH(p[556])) ? `INH(p[556]) : f[596];
        f[597] = 4095;
        f[597] = (f[597] >= `INH(p[558])) ? `INH(p[558]) : f[597];
        f[597] = (f[597] >= `INH(p[559])) ? `INH(p[559]) : f[597];
        f[597] = (f[597] > p[563]) ? p[563] : f[597];
        f[598] = 4095;
        f[598] = (f[598] > p[557]) ? p[557] : f[598];
        f[598] = (f[598] >= `INH(p[563])) ? `INH(p[563]) : f[598];
        f[599] = 4095;
        f[599] = (f[599] > p[561]) ? p[561] : f[599];
        f[599] = (f[599] >= `INH(p[563])) ? `INH(p[563]) : f[599];
        f[600] = 4095;
        f[600] = (f[600] >= p[558]/2) ? p[558]/2 : f[600];
        f[600] = (f[600] >= `INH(p[562])) ? `INH(p[562]) : f[600];
        f[601] = 4095;
        f[601] = (f[601] >= `INH(p[562])) ? `INH(p[562]) : f[601];
        f[601] = (f[601] > p[565]) ? p[565] : f[601];
        f[602] = 4095;
        f[602] = (f[602] > p[558]) ? p[558] : f[602];
        f[602] = (f[602] >= `INH(p[565])) ? `INH(p[565]) : f[602];
        f[602] = (f[602] > p[567]) ? p[567] : f[602];
        f[603] = 4095;
        f[603] = (f[603] >= `INH(p[565])) ? `INH(p[565]) : f[603];
        f[603] = (f[603] > p[568]) ? p[568] : f[603];
        f[604] = 4095;
        f[604] = (f[604] > p[557]) ? p[557] : f[604];
        f[604] = (f[604] >= `INH(p[567])) ? `INH(p[567]) : f[604];
        f[604] = (f[604] >= `INH(p[568])) ? `INH(p[568]) : f[604];
        f[605] = 4095;
        f[605] = (f[605] > p[557]) ? p[557] : f[605];
        f[605] = (f[605] >= `INH(p[566])) ? `INH(p[566]) : f[605];
        f[605] = (f[605] >= `INH(p[568])) ? `INH(p[568]) : f[605];
        f[606] = 4095;
        f[606] = (f[606] >= `INH(p[568])) ? `INH(p[568]) : f[606];
        f[606] = (f[606] > p[570]) ? p[570] : f[606];
        f[607] = 4095;
        f[607] = (f[607] > p[564]) ? p[564] : f[607];
        f[607] = (f[607] >= `INH(p[570])) ? `INH(p[570]) : f[607];
        f[608] = 4095;
        f[608] = (f[608] >= `INH(p[570])) ? `INH(p[570]) : f[608];
        f[608] = (f[608] > p[571]) ? p[571] : f[608];
        f[609] = 4095;
        f[609] = (f[609] > p[569]) ? p[569] : f[609];
        f[609] = (f[609] >= `INH(p[571])) ? `INH(p[571]) : f[609];
        f[610] = 4095;
        f[610] = (f[610] > p[559]) ? p[559] : f[610];
        f[610] = (f[610] > p[566]) ? p[566] : f[610];
        f[610] = (f[610] >= `INH(p[567])) ? `INH(p[567]) : f[610];
        f[610] = (f[610] >= `INH(p[571])) ? `INH(p[571]) : f[610];
        f[611] = 4095;
        f[611] = (f[611] > p[559]) ? p[559] : f[611];
        f[611] = (f[611] >= `INH(p[566])) ? `INH(p[566]) : f[611];
        f[611] = (f[611] >= `INH(p[571])) ? `INH(p[571]) : f[611];
        f[612] = 4095;
        f[612] = (f[612] > p[71]) ? p[71] : f[612];
        f[612] = (f[612] >= `INH(p[573])) ? `INH(p[573]) : f[612];
        f[613] = 4095;
        f[613] = (f[613] > p[572]) ? p[572] : f[613];
        f[613] = (f[613] >= `INH(p[574])) ? `INH(p[574]) : f[613];
        f[614] = 4095;
        f[614] = (f[614] >= `INH(p[71])) ? `INH(p[71]) : f[614];
        f[614] = (f[614] >= `INH(p[573])) ? `INH(p[573]) : f[614];
        f[614] = (f[614] > p[574]) ? p[574] : f[614];
        f[615] = 4095;
        f[615] = (f[615] >= `INH(p[572])) ? `INH(p[572]) : f[615];
        f[615] = (f[615] >= `INH(p[574])) ? `INH(p[574]) : f[615];
        f[615] = (f[615] > p[575]) ? p[575] : f[615];
        f[616] = 4095;
        f[616] = (f[616] > p[72]) ? p[72] : f[616];
        f[616] = (f[616] >= `INH(p[577])) ? `INH(p[577]) : f[616];
        f[617] = 4095;
        f[617] = (f[617] > p[576]) ? p[576] : f[617];
        f[617] = (f[617] >= `INH(p[578])) ? `INH(p[578]) : f[617];
        f[618] = 4095;
        f[618] = (f[618] >= `INH(p[72])) ? `INH(p[72]) : f[618];
        f[618] = (f[618] >= `INH(p[577])) ? `INH(p[577]) : f[618];
        f[618] = (f[618] > p[578]) ? p[578] : f[618];
        f[619] = 4095;
        f[619] = (f[619] >= `INH(p[576])) ? `INH(p[576]) : f[619];
        f[619] = (f[619] >= `INH(p[578])) ? `INH(p[578]) : f[619];
        f[619] = (f[619] > p[579]) ? p[579] : f[619];
        f[620] = 4095;
        f[620] = (f[620] >= `INH(p[21])) ? `INH(p[21]) : f[620];
        f[620] = (f[620] > p[573]) ? p[573] : f[620];
        f[620] = (f[620] > p[577]) ? p[577] : f[620];
        f[621] = 4095;
        f[621] = (f[621] > p[559]) ? p[559] : f[621];
        f[621] = (f[621] >= `INH(p[575])) ? `INH(p[575]) : f[621];
        f[621] = (f[621] >= `INH(p[579])) ? `INH(p[579]) : f[621];
        f[622] = 4095;
        f[622] = (f[622] > p[560]) ? p[560] : f[622];
        f[622] = (f[622] >= `INH(p[580])) ? `INH(p[580]) : f[622];
        f[623] = 4095;
        f[623] = (f[623] > p[73]) ? p[73] : f[623];
        f[623] = (f[623] >= `INH(p[561])) ? `INH(p[561]) : f[623];
        f[624] = 4095;
        f[624] = (f[624] >= `INH(p[73])) ? `INH(p[73]) : f[624];
        f[624] = (f[624] >= `INH(p[561])) ? `INH(p[561]) : f[624];
        f[624] = (f[624] > p[580]) ? p[580] : f[624];
        f[625] = 4095;
        f[625] = (f[625] > p[22]) ? p[22] : f[625];
        f[625] = (f[625] >= `INH(p[560])) ? `INH(p[560]) : f[625];
        f[625] = (f[625] >= `INH(p[580])) ? `INH(p[580]) : f[625];
        f[626] = 4095;
        f[626] = (f[626] >= `INH(p[582])) ? `INH(p[582]) : f[626];
        f[626] = (f[626] >= `INH(p[583])) ? `INH(p[583]) : f[626];
        f[626] = (f[626] > p[587]) ? p[587] : f[626];
        f[627] = 4095;
        f[627] = (f[627] > p[581]) ? p[581] : f[627];
        f[627] = (f[627] >= `INH(p[587])) ? `INH(p[587]) : f[627];
        f[628] = 4095;
        f[628] = (f[628] > p[585]) ? p[585] : f[628];
        f[628] = (f[628] >= `INH(p[587])) ? `INH(p[587]) : f[628];
        f[629] = 4095;
        f[629] = (f[629] >= p[582]/2) ? p[582]/2 : f[629];
        f[629] = (f[629] >= `INH(p[586])) ? `INH(p[586]) : f[629];
        f[630] = 4095;
        f[630] = (f[630] >= `INH(p[586])) ? `INH(p[586]) : f[630];
        f[630] = (f[630] > p[589]) ? p[589] : f[630];
        f[631] = 4095;
        f[631] = (f[631] > p[582]) ? p[582] : f[631];
        f[631] = (f[631] >= `INH(p[589])) ? `INH(p[589]) : f[631];
        f[631] = (f[631] > p[591]) ? p[591] : f[631];
        f[632] = 4095;
        f[632] = (f[632] >= `INH(p[589])) ? `INH(p[589]) : f[632];
        f[632] = (f[632] > p[592]) ? p[592] : f[632];
        f[633] = 4095;
        f[633] = (f[633] > p[581]) ? p[581] : f[633];
        f[633] = (f[633] >= `INH(p[591])) ? `INH(p[591]) : f[633];
        f[633] = (f[633] >= `INH(p[592])) ? `INH(p[592]) : f[633];
        f[634] = 4095;
        f[634] = (f[634] > p[581]) ? p[581] : f[634];
        f[634] = (f[634] >= `INH(p[590])) ? `INH(p[590]) : f[634];
        f[634] = (f[634] >= `INH(p[592])) ? `INH(p[592]) : f[634];
        f[635] = 4095;
        f[635] = (f[635] >= `INH(p[592])) ? `INH(p[592]) : f[635];
        f[635] = (f[635] > p[594]) ? p[594] : f[635];
        f[636] = 4095;
        f[636] = (f[636] > p[588]) ? p[588] : f[636];
        f[636] = (f[636] >= `INH(p[594])) ? `INH(p[594]) : f[636];
        f[637] = 4095;
        f[637] = (f[637] >= `INH(p[594])) ? `INH(p[594]) : f[637];
        f[637] = (f[637] > p[595]) ? p[595] : f[637];
        f[638] = 4095;
        f[638] = (f[638] > p[593]) ? p[593] : f[638];
        f[638] = (f[638] >= `INH(p[595])) ? `INH(p[595]) : f[638];
        f[639] = 4095;
        f[639] = (f[639] > p[583]) ? p[583] : f[639];
        f[639] = (f[639] > p[590]) ? p[590] : f[639];
        f[639] = (f[639] >= `INH(p[591])) ? `INH(p[591]) : f[639];
        f[639] = (f[639] >= `INH(p[595])) ? `INH(p[595]) : f[639];
        f[640] = 4095;
        f[640] = (f[640] > p[583]) ? p[583] : f[640];
        f[640] = (f[640] >= `INH(p[590])) ? `INH(p[590]) : f[640];
        f[640] = (f[640] >= `INH(p[595])) ? `INH(p[595]) : f[640];
        f[641] = 4095;
        f[641] = (f[641] > p[73]) ? p[73] : f[641];
        f[641] = (f[641] >= `INH(p[597])) ? `INH(p[597]) : f[641];
        f[642] = 4095;
        f[642] = (f[642] > p[596]) ? p[596] : f[642];
        f[642] = (f[642] >= `INH(p[598])) ? `INH(p[598]) : f[642];
        f[643] = 4095;
        f[643] = (f[643] >= `INH(p[73])) ? `INH(p[73]) : f[643];
        f[643] = (f[643] >= `INH(p[597])) ? `INH(p[597]) : f[643];
        f[643] = (f[643] > p[598]) ? p[598] : f[643];
        f[644] = 4095;
        f[644] = (f[644] >= `INH(p[596])) ? `INH(p[596]) : f[644];
        f[644] = (f[644] >= `INH(p[598])) ? `INH(p[598]) : f[644];
        f[644] = (f[644] > p[599]) ? p[599] : f[644];
        f[645] = 4095;
        f[645] = (f[645] > p[74]) ? p[74] : f[645];
        f[645] = (f[645] >= `INH(p[601])) ? `INH(p[601]) : f[645];
        f[646] = 4095;
        f[646] = (f[646] > p[600]) ? p[600] : f[646];
        f[646] = (f[646] >= `INH(p[602])) ? `INH(p[602]) : f[646];
        f[647] = 4095;
        f[647] = (f[647] >= `INH(p[74])) ? `INH(p[74]) : f[647];
        f[647] = (f[647] >= `INH(p[601])) ? `INH(p[601]) : f[647];
        f[647] = (f[647] > p[602]) ? p[602] : f[647];
        f[648] = 4095;
        f[648] = (f[648] >= `INH(p[600])) ? `INH(p[600]) : f[648];
        f[648] = (f[648] >= `INH(p[602])) ? `INH(p[602]) : f[648];
        f[648] = (f[648] > p[603]) ? p[603] : f[648];
        f[649] = 4095;
        f[649] = (f[649] >= `INH(p[22])) ? `INH(p[22]) : f[649];
        f[649] = (f[649] > p[597]) ? p[597] : f[649];
        f[649] = (f[649] > p[601]) ? p[601] : f[649];
        f[650] = 4095;
        f[650] = (f[650] > p[583]) ? p[583] : f[650];
        f[650] = (f[650] >= `INH(p[599])) ? `INH(p[599]) : f[650];
        f[650] = (f[650] >= `INH(p[603])) ? `INH(p[603]) : f[650];
        f[651] = 4095;
        f[651] = (f[651] > p[584]) ? p[584] : f[651];
        f[651] = (f[651] >= `INH(p[604])) ? `INH(p[604]) : f[651];
        f[652] = 4095;
        f[652] = (f[652] > p[75]) ? p[75] : f[652];
        f[652] = (f[652] >= `INH(p[585])) ? `INH(p[585]) : f[652];
        f[653] = 4095;
        f[653] = (f[653] >= `INH(p[75])) ? `INH(p[75]) : f[653];
        f[653] = (f[653] >= `INH(p[585])) ? `INH(p[585]) : f[653];
        f[653] = (f[653] > p[604]) ? p[604] : f[653];
        f[654] = 4095;
        f[654] = (f[654] > p[23]) ? p[23] : f[654];
        f[654] = (f[654] >= `INH(p[584])) ? `INH(p[584]) : f[654];
        f[654] = (f[654] >= `INH(p[604])) ? `INH(p[604]) : f[654];
        f[655] = 4095;
        f[655] = (f[655] > p[606]) ? p[606] : f[655];
        f[655] = (f[655] >= `INH(p[608])) ? `INH(p[608]) : f[655];
        f[656] = 4095;
        f[656] = (f[656] >= `INH(p[605])) ? `INH(p[605]) : f[656];
        f[656] = (f[656] >= `INH(p[606])) ? `INH(p[606]) : f[656];
        f[656] = (f[656] >= `INH(p[608])) ? `INH(p[608]) : f[656];
        f[656] = (f[656] > p[609]) ? p[609] : f[656];
        f[657] = 4095;
        f[657] = (f[657] > p[75]) ? p[75] : f[657];
        f[657] = (f[657] >= `INH(p[611])) ? `INH(p[611]) : f[657];
        f[658] = 4095;
        f[658] = (f[658] > p[610]) ? p[610] : f[658];
        f[658] = (f[658] >= `INH(p[612])) ? `INH(p[612]) : f[658];
        f[659] = 4095;
        f[659] = (f[659] >= `INH(p[75])) ? `INH(p[75]) : f[659];
        f[659] = (f[659] >= `INH(p[611])) ? `INH(p[611]) : f[659];
        f[659] = (f[659] > p[612]) ? p[612] : f[659];
        f[660] = 4095;
        f[660] = (f[660] >= `INH(p[610])) ? `INH(p[610]) : f[660];
        f[660] = (f[660] >= `INH(p[612])) ? `INH(p[612]) : f[660];
        f[660] = (f[660] > p[613]) ? p[613] : f[660];
        f[661] = 4095;
        f[661] = (f[661] > p[70]) ? p[70] : f[661];
        f[661] = (f[661] >= `INH(p[615])) ? `INH(p[615]) : f[661];
        f[662] = 4095;
        f[662] = (f[662] > p[614]) ? p[614] : f[662];
        f[662] = (f[662] >= `INH(p[616])) ? `INH(p[616]) : f[662];
        f[663] = 4095;
        f[663] = (f[663] >= `INH(p[70])) ? `INH(p[70]) : f[663];
        f[663] = (f[663] >= `INH(p[615])) ? `INH(p[615]) : f[663];
        f[663] = (f[663] > p[616]) ? p[616] : f[663];
        f[664] = 4095;
        f[664] = (f[664] >= `INH(p[614])) ? `INH(p[614]) : f[664];
        f[664] = (f[664] >= `INH(p[616])) ? `INH(p[616]) : f[664];
        f[664] = (f[664] > p[617]) ? p[617] : f[664];
        f[665] = 4095;
        f[665] = (f[665] >= `INH(p[23])) ? `INH(p[23]) : f[665];
        f[665] = (f[665] > p[611]) ? p[611] : f[665];
        f[665] = (f[665] > p[615]) ? p[615] : f[665];
        f[666] = 4095;
        f[666] = (f[666] > p[608]) ? p[608] : f[666];
        f[666] = (f[666] >= `INH(p[613])) ? `INH(p[613]) : f[666];
        f[666] = (f[666] >= `INH(p[617])) ? `INH(p[617]) : f[666];
        f[667] = 4095;
        f[667] = (f[667] > p[607]) ? p[607] : f[667];
        f[667] = (f[667] >= `INH(p[618])) ? `INH(p[618]) : f[667];
        f[668] = 4095;
        f[668] = (f[668] > p[76]) ? p[76] : f[668];
        f[668] = (f[668] >= `INH(p[609])) ? `INH(p[609]) : f[668];
        f[669] = 4095;
        f[669] = (f[669] >= `INH(p[76])) ? `INH(p[76]) : f[669];
        f[669] = (f[669] >= `INH(p[609])) ? `INH(p[609]) : f[669];
        f[669] = (f[669] > p[618]) ? p[618] : f[669];
        f[670] = 4095;
        f[670] = (f[670] > p[24]) ? p[24] : f[670];
        f[670] = (f[670] >= `INH(p[607])) ? `INH(p[607]) : f[670];
        f[670] = (f[670] >= `INH(p[618])) ? `INH(p[618]) : f[670];
        f[671] = 4095;
        f[671] = (f[671] >= `INH(p[620])) ? `INH(p[620]) : f[671];
        f[671] = (f[671] >= `INH(p[621])) ? `INH(p[621]) : f[671];
        f[671] = (f[671] > p[625]) ? p[625] : f[671];
        f[672] = 4095;
        f[672] = (f[672] > p[619]) ? p[619] : f[672];
        f[672] = (f[672] >= `INH(p[625])) ? `INH(p[625]) : f[672];
        f[673] = 4095;
        f[673] = (f[673] > p[623]) ? p[623] : f[673];
        f[673] = (f[673] >= `INH(p[625])) ? `INH(p[625]) : f[673];
        f[674] = 4095;
        f[674] = (f[674] >= p[620]/2) ? p[620]/2 : f[674];
        f[674] = (f[674] >= `INH(p[624])) ? `INH(p[624]) : f[674];
        f[675] = 4095;
        f[675] = (f[675] >= `INH(p[624])) ? `INH(p[624]) : f[675];
        f[675] = (f[675] > p[627]) ? p[627] : f[675];
        f[676] = 4095;
        f[676] = (f[676] > p[620]) ? p[620] : f[676];
        f[676] = (f[676] >= `INH(p[627])) ? `INH(p[627]) : f[676];
        f[676] = (f[676] > p[629]) ? p[629] : f[676];
        f[677] = 4095;
        f[677] = (f[677] >= `INH(p[627])) ? `INH(p[627]) : f[677];
        f[677] = (f[677] > p[630]) ? p[630] : f[677];
        f[678] = 4095;
        f[678] = (f[678] > p[619]) ? p[619] : f[678];
        f[678] = (f[678] >= `INH(p[629])) ? `INH(p[629]) : f[678];
        f[678] = (f[678] >= `INH(p[630])) ? `INH(p[630]) : f[678];
        f[679] = 4095;
        f[679] = (f[679] > p[619]) ? p[619] : f[679];
        f[679] = (f[679] >= `INH(p[628])) ? `INH(p[628]) : f[679];
        f[679] = (f[679] >= `INH(p[630])) ? `INH(p[630]) : f[679];
        f[680] = 4095;
        f[680] = (f[680] >= `INH(p[630])) ? `INH(p[630]) : f[680];
        f[680] = (f[680] > p[632]) ? p[632] : f[680];
        f[681] = 4095;
        f[681] = (f[681] > p[626]) ? p[626] : f[681];
        f[681] = (f[681] >= `INH(p[632])) ? `INH(p[632]) : f[681];
        f[682] = 4095;
        f[682] = (f[682] >= `INH(p[632])) ? `INH(p[632]) : f[682];
        f[682] = (f[682] > p[633]) ? p[633] : f[682];
        f[683] = 4095;
        f[683] = (f[683] > p[631]) ? p[631] : f[683];
        f[683] = (f[683] >= `INH(p[633])) ? `INH(p[633]) : f[683];
        f[684] = 4095;
        f[684] = (f[684] > p[621]) ? p[621] : f[684];
        f[684] = (f[684] > p[628]) ? p[628] : f[684];
        f[684] = (f[684] >= `INH(p[629])) ? `INH(p[629]) : f[684];
        f[684] = (f[684] >= `INH(p[633])) ? `INH(p[633]) : f[684];
        f[685] = 4095;
        f[685] = (f[685] > p[621]) ? p[621] : f[685];
        f[685] = (f[685] >= `INH(p[628])) ? `INH(p[628]) : f[685];
        f[685] = (f[685] >= `INH(p[633])) ? `INH(p[633]) : f[685];
        f[686] = 4095;
        f[686] = (f[686] > p[77]) ? p[77] : f[686];
        f[686] = (f[686] >= `INH(p[635])) ? `INH(p[635]) : f[686];
        f[687] = 4095;
        f[687] = (f[687] > p[634]) ? p[634] : f[687];
        f[687] = (f[687] >= `INH(p[636])) ? `INH(p[636]) : f[687];
        f[688] = 4095;
        f[688] = (f[688] >= `INH(p[77])) ? `INH(p[77]) : f[688];
        f[688] = (f[688] >= `INH(p[635])) ? `INH(p[635]) : f[688];
        f[688] = (f[688] > p[636]) ? p[636] : f[688];
        f[689] = 4095;
        f[689] = (f[689] >= `INH(p[634])) ? `INH(p[634]) : f[689];
        f[689] = (f[689] >= `INH(p[636])) ? `INH(p[636]) : f[689];
        f[689] = (f[689] > p[637]) ? p[637] : f[689];
        f[690] = 4095;
        f[690] = (f[690] > p[78]) ? p[78] : f[690];
        f[690] = (f[690] >= `INH(p[639])) ? `INH(p[639]) : f[690];
        f[691] = 4095;
        f[691] = (f[691] > p[638]) ? p[638] : f[691];
        f[691] = (f[691] >= `INH(p[640])) ? `INH(p[640]) : f[691];
        f[692] = 4095;
        f[692] = (f[692] >= `INH(p[78])) ? `INH(p[78]) : f[692];
        f[692] = (f[692] >= `INH(p[639])) ? `INH(p[639]) : f[692];
        f[692] = (f[692] > p[640]) ? p[640] : f[692];
        f[693] = 4095;
        f[693] = (f[693] >= `INH(p[638])) ? `INH(p[638]) : f[693];
        f[693] = (f[693] >= `INH(p[640])) ? `INH(p[640]) : f[693];
        f[693] = (f[693] > p[641]) ? p[641] : f[693];
        f[694] = 4095;
        f[694] = (f[694] >= `INH(p[24])) ? `INH(p[24]) : f[694];
        f[694] = (f[694] > p[635]) ? p[635] : f[694];
        f[694] = (f[694] > p[639]) ? p[639] : f[694];
        f[695] = 4095;
        f[695] = (f[695] > p[621]) ? p[621] : f[695];
        f[695] = (f[695] >= `INH(p[637])) ? `INH(p[637]) : f[695];
        f[695] = (f[695] >= `INH(p[641])) ? `INH(p[641]) : f[695];
        f[696] = 4095;
        f[696] = (f[696] > p[622]) ? p[622] : f[696];
        f[696] = (f[696] >= `INH(p[642])) ? `INH(p[642]) : f[696];
        f[697] = 4095;
        f[697] = (f[697] > p[79]) ? p[79] : f[697];
        f[697] = (f[697] >= `INH(p[623])) ? `INH(p[623]) : f[697];
        f[698] = 4095;
        f[698] = (f[698] >= `INH(p[79])) ? `INH(p[79]) : f[698];
        f[698] = (f[698] >= `INH(p[623])) ? `INH(p[623]) : f[698];
        f[698] = (f[698] > p[642]) ? p[642] : f[698];
        f[699] = 4095;
        f[699] = (f[699] > p[25]) ? p[25] : f[699];
        f[699] = (f[699] >= `INH(p[622])) ? `INH(p[622]) : f[699];
        f[699] = (f[699] >= `INH(p[642])) ? `INH(p[642]) : f[699];
        f[700] = 4095;
        f[700] = (f[700] > p[644]) ? p[644] : f[700];
        f[700] = (f[700] >= `INH(p[646])) ? `INH(p[646]) : f[700];
        f[701] = 4095;
        f[701] = (f[701] >= `INH(p[643])) ? `INH(p[643]) : f[701];
        f[701] = (f[701] >= `INH(p[644])) ? `INH(p[644]) : f[701];
        f[701] = (f[701] >= `INH(p[646])) ? `INH(p[646]) : f[701];
        f[701] = (f[701] > p[647]) ? p[647] : f[701];
        f[702] = 4095;
        f[702] = (f[702] > p[79]) ? p[79] : f[702];
        f[702] = (f[702] >= `INH(p[649])) ? `INH(p[649]) : f[702];
        f[703] = 4095;
        f[703] = (f[703] > p[648]) ? p[648] : f[703];
        f[703] = (f[703] >= `INH(p[650])) ? `INH(p[650]) : f[703];
        f[704] = 4095;
        f[704] = (f[704] >= `INH(p[79])) ? `INH(p[79]) : f[704];
        f[704] = (f[704] >= `INH(p[649])) ? `INH(p[649]) : f[704];
        f[704] = (f[704] > p[650]) ? p[650] : f[704];
        f[705] = 4095;
        f[705] = (f[705] >= `INH(p[648])) ? `INH(p[648]) : f[705];
        f[705] = (f[705] >= `INH(p[650])) ? `INH(p[650]) : f[705];
        f[705] = (f[705] > p[651]) ? p[651] : f[705];
        f[706] = 4095;
        f[706] = (f[706] > p[76]) ? p[76] : f[706];
        f[706] = (f[706] >= `INH(p[653])) ? `INH(p[653]) : f[706];
        f[707] = 4095;
        f[707] = (f[707] > p[652]) ? p[652] : f[707];
        f[707] = (f[707] >= `INH(p[654])) ? `INH(p[654]) : f[707];
        f[708] = 4095;
        f[708] = (f[708] >= `INH(p[76])) ? `INH(p[76]) : f[708];
        f[708] = (f[708] >= `INH(p[653])) ? `INH(p[653]) : f[708];
        f[708] = (f[708] > p[654]) ? p[654] : f[708];
        f[709] = 4095;
        f[709] = (f[709] >= `INH(p[652])) ? `INH(p[652]) : f[709];
        f[709] = (f[709] >= `INH(p[654])) ? `INH(p[654]) : f[709];
        f[709] = (f[709] > p[655]) ? p[655] : f[709];
        f[710] = 4095;
        f[710] = (f[710] >= `INH(p[25])) ? `INH(p[25]) : f[710];
        f[710] = (f[710] > p[649]) ? p[649] : f[710];
        f[710] = (f[710] > p[653]) ? p[653] : f[710];
        f[711] = 4095;
        f[711] = (f[711] > p[646]) ? p[646] : f[711];
        f[711] = (f[711] >= `INH(p[651])) ? `INH(p[651]) : f[711];
        f[711] = (f[711] >= `INH(p[655])) ? `INH(p[655]) : f[711];
        f[712] = 4095;
        f[712] = (f[712] > p[645]) ? p[645] : f[712];
        f[712] = (f[712] >= `INH(p[656])) ? `INH(p[656]) : f[712];
        f[713] = 4095;
        f[713] = (f[713] > p[80]) ? p[80] : f[713];
        f[713] = (f[713] >= `INH(p[647])) ? `INH(p[647]) : f[713];
        f[714] = 4095;
        f[714] = (f[714] >= `INH(p[80])) ? `INH(p[80]) : f[714];
        f[714] = (f[714] >= `INH(p[647])) ? `INH(p[647]) : f[714];
        f[714] = (f[714] > p[656]) ? p[656] : f[714];
        f[715] = 4095;
        f[715] = (f[715] > p[26]) ? p[26] : f[715];
        f[715] = (f[715] >= `INH(p[645])) ? `INH(p[645]) : f[715];
        f[715] = (f[715] >= `INH(p[656])) ? `INH(p[656]) : f[715];
        f[716] = 4095;
        f[716] = (f[716] > p[658]) ? p[658] : f[716];
        f[716] = (f[716] >= `INH(p[660])) ? `INH(p[660]) : f[716];
        f[717] = 4095;
        f[717] = (f[717] >= `INH(p[657])) ? `INH(p[657]) : f[717];
        f[717] = (f[717] >= `INH(p[658])) ? `INH(p[658]) : f[717];
        f[717] = (f[717] >= `INH(p[660])) ? `INH(p[660]) : f[717];
        f[717] = (f[717] > p[661]) ? p[661] : f[717];
        f[718] = 4095;
        f[718] = (f[718] > p[80]) ? p[80] : f[718];
        f[718] = (f[718] >= `INH(p[663])) ? `INH(p[663]) : f[718];
        f[719] = 4095;
        f[719] = (f[719] > p[662]) ? p[662] : f[719];
        f[719] = (f[719] >= `INH(p[664])) ? `INH(p[664]) : f[719];
        f[720] = 4095;
        f[720] = (f[720] >= `INH(p[80])) ? `INH(p[80]) : f[720];
        f[720] = (f[720] >= `INH(p[663])) ? `INH(p[663]) : f[720];
        f[720] = (f[720] > p[664]) ? p[664] : f[720];
        f[721] = 4095;
        f[721] = (f[721] >= `INH(p[662])) ? `INH(p[662]) : f[721];
        f[721] = (f[721] >= `INH(p[664])) ? `INH(p[664]) : f[721];
        f[721] = (f[721] > p[665]) ? p[665] : f[721];
        f[722] = 4095;
        f[722] = (f[722] > p[81]) ? p[81] : f[722];
        f[722] = (f[722] >= `INH(p[667])) ? `INH(p[667]) : f[722];
        f[723] = 4095;
        f[723] = (f[723] > p[666]) ? p[666] : f[723];
        f[723] = (f[723] >= `INH(p[668])) ? `INH(p[668]) : f[723];
        f[724] = 4095;
        f[724] = (f[724] >= `INH(p[81])) ? `INH(p[81]) : f[724];
        f[724] = (f[724] >= `INH(p[667])) ? `INH(p[667]) : f[724];
        f[724] = (f[724] > p[668]) ? p[668] : f[724];
        f[725] = 4095;
        f[725] = (f[725] >= `INH(p[666])) ? `INH(p[666]) : f[725];
        f[725] = (f[725] >= `INH(p[668])) ? `INH(p[668]) : f[725];
        f[725] = (f[725] > p[669]) ? p[669] : f[725];
        f[726] = 4095;
        f[726] = (f[726] >= `INH(p[26])) ? `INH(p[26]) : f[726];
        f[726] = (f[726] > p[663]) ? p[663] : f[726];
        f[726] = (f[726] > p[667]) ? p[667] : f[726];
        f[727] = 4095;
        f[727] = (f[727] > p[660]) ? p[660] : f[727];
        f[727] = (f[727] >= `INH(p[665])) ? `INH(p[665]) : f[727];
        f[727] = (f[727] >= `INH(p[669])) ? `INH(p[669]) : f[727];
        f[728] = 4095;
        f[728] = (f[728] > p[659]) ? p[659] : f[728];
        f[728] = (f[728] >= `INH(p[670])) ? `INH(p[670]) : f[728];
        f[729] = 4095;
        f[729] = (f[729] > p[82]) ? p[82] : f[729];
        f[729] = (f[729] >= `INH(p[661])) ? `INH(p[661]) : f[729];
        f[730] = 4095;
        f[730] = (f[730] >= `INH(p[82])) ? `INH(p[82]) : f[730];
        f[730] = (f[730] >= `INH(p[661])) ? `INH(p[661]) : f[730];
        f[730] = (f[730] > p[670]) ? p[670] : f[730];
        f[731] = 4095;
        f[731] = (f[731] > p[27]) ? p[27] : f[731];
        f[731] = (f[731] >= `INH(p[659])) ? `INH(p[659]) : f[731];
        f[731] = (f[731] >= `INH(p[670])) ? `INH(p[670]) : f[731];
        if(f[27]>0)
                f[0] = 0;
        if(f[28]>0)
                f[29] = 0;
        if(f[30]>0)
                f[31] = 0;
        if(f[32]>0)
                f[33] = 0;
        if(f[34]>0)
                f[36] = 0;
        if(f[35]>0)
                f[36] = 0;
        if(f[37]>0)
                f[38] = 0;
        if(f[39]>0)
                f[40] = 0;
        if(f[39]>0)
                f[41] = 0;
        if(f[56]>0)
                f[1] = 0;
        if(f[57]>0)
                f[58] = 0;
        if(f[59]>0)
                f[60] = 0;
        if(f[61]>0)
                f[62] = 0;
        if(f[63]>0)
                f[65] = 0;
        if(f[64]>0)
                f[65] = 0;
        if(f[66]>0)
                f[67] = 0;
        if(f[68]>0)
                f[69] = 0;
        if(f[68]>0)
                f[70] = 0;
        if(f[85]>0)
                f[2] = 0;
        if(f[86]>0)
                f[87] = 0;
        if(f[88]>0)
                f[89] = 0;
        if(f[90]>0)
                f[91] = 0;
        if(f[92]>0)
                f[94] = 0;
        if(f[93]>0)
                f[94] = 0;
        if(f[95]>0)
                f[96] = 0;
        if(f[97]>0)
                f[98] = 0;
        if(f[97]>0)
                f[99] = 0;
        if(f[114]>0)
                f[3] = 0;
        if(f[115]>0)
                f[116] = 0;
        if(f[117]>0)
                f[118] = 0;
        if(f[119]>0)
                f[120] = 0;
        if(f[121]>0)
                f[123] = 0;
        if(f[122]>0)
                f[123] = 0;
        if(f[124]>0)
                f[125] = 0;
        if(f[126]>0)
                f[127] = 0;
        if(f[126]>0)
                f[128] = 0;
        if(f[143]>0)
                f[4] = 0;
        if(f[144]>0)
                f[145] = 0;
        if(f[146]>0)
                f[147] = 0;
        if(f[148]>0)
                f[149] = 0;
        if(f[150]>0)
                f[152] = 0;
        if(f[151]>0)
                f[152] = 0;
        if(f[153]>0)
                f[154] = 0;
        if(f[155]>0)
                f[156] = 0;
        if(f[155]>0)
                f[157] = 0;
        if(f[172]>0)
                f[5] = 0;
        if(f[173]>0)
                f[174] = 0;
        if(f[175]>0)
                f[176] = 0;
        if(f[177]>0)
                f[178] = 0;
        if(f[179]>0)
                f[181] = 0;
        if(f[180]>0)
                f[181] = 0;
        if(f[182]>0)
                f[183] = 0;
        if(f[184]>0)
                f[185] = 0;
        if(f[184]>0)
                f[186] = 0;
        if(f[201]>0)
                f[6] = 0;
        if(f[202]>0)
                f[203] = 0;
        if(f[204]>0)
                f[205] = 0;
        if(f[206]>0)
                f[207] = 0;
        if(f[208]>0)
                f[210] = 0;
        if(f[209]>0)
                f[210] = 0;
        if(f[211]>0)
                f[212] = 0;
        if(f[213]>0)
                f[214] = 0;
        if(f[213]>0)
                f[215] = 0;
        if(f[230]>0)
                f[7] = 0;
        if(f[231]>0)
                f[232] = 0;
        if(f[233]>0)
                f[234] = 0;
        if(f[235]>0)
                f[236] = 0;
        if(f[237]>0)
                f[239] = 0;
        if(f[238]>0)
                f[239] = 0;
        if(f[240]>0)
                f[241] = 0;
        if(f[242]>0)
                f[243] = 0;
        if(f[242]>0)
                f[244] = 0;
        if(f[259]>0)
                f[8] = 0;
        if(f[260]>0)
                f[261] = 0;
        if(f[262]>0)
                f[263] = 0;
        if(f[264]>0)
                f[265] = 0;
        if(f[266]>0)
                f[268] = 0;
        if(f[267]>0)
                f[268] = 0;
        if(f[269]>0)
                f[270] = 0;
        if(f[271]>0)
                f[272] = 0;
        if(f[271]>0)
                f[273] = 0;
        if(f[288]>0)
                f[9] = 0;
        if(f[289]>0)
                f[290] = 0;
        if(f[291]>0)
                f[292] = 0;
        if(f[293]>0)
                f[294] = 0;
        if(f[295]>0)
                f[297] = 0;
        if(f[296]>0)
                f[297] = 0;
        if(f[298]>0)
                f[299] = 0;
        if(f[300]>0)
                f[301] = 0;
        if(f[300]>0)
                f[302] = 0;
        if(f[317]>0)
                f[10] = 0;
        if(f[318]>0)
                f[319] = 0;
        if(f[320]>0)
                f[321] = 0;
        if(f[322]>0)
                f[323] = 0;
        if(f[324]>0)
                f[326] = 0;
        if(f[325]>0)
                f[326] = 0;
        if(f[327]>0)
                f[328] = 0;
        if(f[329]>0)
                f[330] = 0;
        if(f[329]>0)
                f[331] = 0;
        if(f[362]>0)
                f[12] = 0;
        if(f[363]>0)
                f[364] = 0;
        if(f[365]>0)
                f[366] = 0;
        if(f[367]>0)
                f[368] = 0;
        if(f[369]>0)
                f[371] = 0;
        if(f[370]>0)
                f[371] = 0;
        if(f[372]>0)
                f[373] = 0;
        if(f[374]>0)
                f[375] = 0;
        if(f[374]>0)
                f[376] = 0;
        if(f[391]>0)
                f[13] = 0;
        if(f[392]>0)
                f[393] = 0;
        if(f[394]>0)
                f[395] = 0;
        if(f[396]>0)
                f[397] = 0;
        if(f[398]>0)
                f[400] = 0;
        if(f[399]>0)
                f[400] = 0;
        if(f[401]>0)
                f[402] = 0;
        if(f[403]>0)
                f[404] = 0;
        if(f[403]>0)
                f[405] = 0;
        if(f[420]>0)
                f[14] = 0;
        if(f[421]>0)
                f[422] = 0;
        if(f[423]>0)
                f[424] = 0;
        if(f[425]>0)
                f[426] = 0;
        if(f[427]>0)
                f[429] = 0;
        if(f[428]>0)
                f[429] = 0;
        if(f[430]>0)
                f[431] = 0;
        if(f[432]>0)
                f[433] = 0;
        if(f[432]>0)
                f[434] = 0;
        if(f[449]>0)
                f[15] = 0;
        if(f[450]>0)
                f[451] = 0;
        if(f[452]>0)
                f[453] = 0;
        if(f[454]>0)
                f[455] = 0;
        if(f[456]>0)
                f[458] = 0;
        if(f[457]>0)
                f[458] = 0;
        if(f[459]>0)
                f[460] = 0;
        if(f[461]>0)
                f[462] = 0;
        if(f[461]>0)
                f[463] = 0;
        if(f[494]>0)
                f[17] = 0;
        if(f[495]>0)
                f[496] = 0;
        if(f[497]>0)
                f[498] = 0;
        if(f[499]>0)
                f[500] = 0;
        if(f[501]>0)
                f[503] = 0;
        if(f[502]>0)
                f[503] = 0;
        if(f[504]>0)
                f[505] = 0;
        if(f[506]>0)
                f[507] = 0;
        if(f[506]>0)
                f[508] = 0;
        if(f[523]>0)
                f[18] = 0;
        if(f[524]>0)
                f[525] = 0;
        if(f[526]>0)
                f[527] = 0;
        if(f[528]>0)
                f[529] = 0;
        if(f[530]>0)
                f[532] = 0;
        if(f[531]>0)
                f[532] = 0;
        if(f[533]>0)
                f[534] = 0;
        if(f[535]>0)
                f[536] = 0;
        if(f[535]>0)
                f[537] = 0;
        if(f[552]>0)
                f[19] = 0;
        if(f[553]>0)
                f[554] = 0;
        if(f[555]>0)
                f[556] = 0;
        if(f[557]>0)
                f[558] = 0;
        if(f[559]>0)
                f[561] = 0;
        if(f[560]>0)
                f[561] = 0;
        if(f[562]>0)
                f[563] = 0;
        if(f[564]>0)
                f[565] = 0;
        if(f[564]>0)
                f[566] = 0;
        if(f[597]>0)
                f[21] = 0;
        if(f[598]>0)
                f[599] = 0;
        if(f[600]>0)
                f[601] = 0;
        if(f[602]>0)
                f[603] = 0;
        if(f[604]>0)
                f[606] = 0;
        if(f[605]>0)
                f[606] = 0;
        if(f[607]>0)
                f[608] = 0;
        if(f[609]>0)
                f[610] = 0;
        if(f[609]>0)
                f[611] = 0;
        if(f[626]>0)
                f[22] = 0;
        if(f[627]>0)
                f[628] = 0;
        if(f[629]>0)
                f[630] = 0;
        if(f[631]>0)
                f[632] = 0;
        if(f[633]>0)
                f[635] = 0;
        if(f[634]>0)
                f[635] = 0;
        if(f[636]>0)
                f[637] = 0;
        if(f[638]>0)
                f[639] = 0;
        if(f[638]>0)
                f[640] = 0;
        if(f[671]>0)
                f[24] = 0;
        if(f[672]>0)
                f[673] = 0;
        if(f[674]>0)
                f[675] = 0;
        if(f[676]>0)
                f[677] = 0;
        if(f[678]>0)
                f[680] = 0;
        if(f[679]>0)
                f[680] = 0;
        if(f[681]>0)
                f[682] = 0;
        if(f[683]>0)
                f[684] = 0;
        if(f[683]>0)
                f[685] = 0;
        tf = (f[0]>0)?1:(f[1]>0)?2:(f[2]>0)?3:(f[3]>0)?4:(f[4]>0)?5:(f[5]>0)?6:(f[6]>0)?7:(f[7]>0)?8:(f[8]>0)?9:(f[9]>0)?10:(f[10]>0)?11:(f[11]>0)?12:(f[12]>0)?13:(f[13]>0)?14:(f[14]>0)?15:(f[15]>0)?16:(f[16]>0)?17:(f[17]>0)?18:(f[18]>0)?19:(f[19]>0)?20:(f[20]>0)?21:(f[21]>0)?22:(f[22]>0)?23:(f[23]>0)?24:(f[24]>0)?25:(f[25]>0)?26:(f[26]>0)?27:(f[27]>0)?28:(f[28]>0)?29:(f[29]>0)?30:(f[30]>0)?31:(f[31]>0)?32:(f[32]>0)?33:(f[33]>0)?34:(f[34]>0)?35:(f[35]>0)?36:(f[36]>0)?37:(f[37]>0)?38:(f[38]>0)?39:(f[39]>0)?40:(f[40]>0)?41:(f[41]>0)?42:(f[42]>0)?43:(f[43]>0)?44:(f[44]>0)?45:(f[45]>0)?46:(f[46]>0)?47:(f[47]>0)?48:(f[48]>0)?49:(f[49]>0)?50:(f[50]>0)?51:(f[51]>0)?52:(f[52]>0)?53:(f[53]>0)?54:(f[54]>0)?55:(f[55]>0)?56:(f[56]>0)?57:(f[57]>0)?58:(f[58]>0)?59:(f[59]>0)?60:(f[60]>0)?61:(f[61]>0)?62:(f[62]>0)?63:(f[63]>0)?64:(f[64]>0)?65:(f[65]>0)?66:(f[66]>0)?67:(f[67]>0)?68:(f[68]>0)?69:(f[69]>0)?70:(f[70]>0)?71:(f[71]>0)?72:(f[72]>0)?73:(f[73]>0)?74:(f[74]>0)?75:(f[75]>0)?76:(f[76]>0)?77:(f[77]>0)?78:(f[78]>0)?79:(f[79]>0)?80:(f[80]>0)?81:(f[81]>0)?82:(f[82]>0)?83:(f[83]>0)?84:(f[84]>0)?85:(f[85]>0)?86:(f[86]>0)?87:(f[87]>0)?88:(f[88]>0)?89:(f[89]>0)?90:(f[90]>0)?91:(f[91]>0)?92:(f[92]>0)?93:(f[93]>0)?94:(f[94]>0)?95:(f[95]>0)?96:(f[96]>0)?97:(f[97]>0)?98:(f[98]>0)?99:(f[99]>0)?100:(f[100]>0)?101:(f[101]>0)?102:(f[102]>0)?103:(f[103]>0)?104:(f[104]>0)?105:(f[105]>0)?106:(f[106]>0)?107:(f[107]>0)?108:(f[108]>0)?109:(f[109]>0)?110:(f[110]>0)?111:(f[111]>0)?112:(f[112]>0)?113:(f[113]>0)?114:(f[114]>0)?115:(f[115]>0)?116:(f[116]>0)?117:(f[117]>0)?118:(f[118]>0)?119:(f[119]>0)?120:(f[120]>0)?121:(f[121]>0)?122:(f[122]>0)?123:(f[123]>0)?124:(f[124]>0)?125:(f[125]>0)?126:(f[126]>0)?127:(f[127]>0)?128:(f[128]>0)?129:(f[129]>0)?130:(f[130]>0)?131:(f[131]>0)?132:(f[132]>0)?133:(f[133]>0)?134:(f[134]>0)?135:(f[135]>0)?136:(f[136]>0)?137:(f[137]>0)?138:(f[138]>0)?139:(f[139]>0)?140:(f[140]>0)?141:(f[141]>0)?142:(f[142]>0)?143:(f[143]>0)?144:(f[144]>0)?145:(f[145]>0)?146:(f[146]>0)?147:(f[147]>0)?148:(f[148]>0)?149:(f[149]>0)?150:(f[150]>0)?151:(f[151]>0)?152:(f[152]>0)?153:(f[153]>0)?154:(f[154]>0)?155:(f[155]>0)?156:(f[156]>0)?157:(f[157]>0)?158:(f[158]>0)?159:(f[159]>0)?160:(f[160]>0)?161:(f[161]>0)?162:(f[162]>0)?163:(f[163]>0)?164:(f[164]>0)?165:(f[165]>0)?166:(f[166]>0)?167:(f[167]>0)?168:(f[168]>0)?169:(f[169]>0)?170:(f[170]>0)?171:(f[171]>0)?172:(f[172]>0)?173:(f[173]>0)?174:(f[174]>0)?175:(f[175]>0)?176:(f[176]>0)?177:(f[177]>0)?178:(f[178]>0)?179:(f[179]>0)?180:(f[180]>0)?181:(f[181]>0)?182:(f[182]>0)?183:(f[183]>0)?184:(f[184]>0)?185:(f[185]>0)?186:(f[186]>0)?187:(f[187]>0)?188:(f[188]>0)?189:(f[189]>0)?190:(f[190]>0)?191:(f[191]>0)?192:(f[192]>0)?193:(f[193]>0)?194:(f[194]>0)?195:(f[195]>0)?196:(f[196]>0)?197:(f[197]>0)?198:(f[198]>0)?199:(f[199]>0)?200:(f[200]>0)?201:(f[201]>0)?202:(f[202]>0)?203:(f[203]>0)?204:(f[204]>0)?205:(f[205]>0)?206:(f[206]>0)?207:(f[207]>0)?208:(f[208]>0)?209:(f[209]>0)?210:(f[210]>0)?211:(f[211]>0)?212:(f[212]>0)?213:(f[213]>0)?214:(f[214]>0)?215:(f[215]>0)?216:(f[216]>0)?217:(f[217]>0)?218:(f[218]>0)?219:(f[219]>0)?220:(f[220]>0)?221:(f[221]>0)?222:(f[222]>0)?223:(f[223]>0)?224:(f[224]>0)?225:(f[225]>0)?226:(f[226]>0)?227:(f[227]>0)?228:(f[228]>0)?229:(f[229]>0)?230:(f[230]>0)?231:(f[231]>0)?232:(f[232]>0)?233:(f[233]>0)?234:(f[234]>0)?235:(f[235]>0)?236:(f[236]>0)?237:(f[237]>0)?238:(f[238]>0)?239:(f[239]>0)?240:(f[240]>0)?241:(f[241]>0)?242:(f[242]>0)?243:(f[243]>0)?244:(f[244]>0)?245:(f[245]>0)?246:(f[246]>0)?247:(f[247]>0)?248:(f[248]>0)?249:(f[249]>0)?250:(f[250]>0)?251:(f[251]>0)?252:(f[252]>0)?253:(f[253]>0)?254:(f[254]>0)?255:(f[255]>0)?256:(f[256]>0)?257:(f[257]>0)?258:(f[258]>0)?259:(f[259]>0)?260:(f[260]>0)?261:(f[261]>0)?262:(f[262]>0)?263:(f[263]>0)?264:(f[264]>0)?265:(f[265]>0)?266:(f[266]>0)?267:(f[267]>0)?268:(f[268]>0)?269:(f[269]>0)?270:(f[270]>0)?271:(f[271]>0)?272:(f[272]>0)?273:(f[273]>0)?274:(f[274]>0)?275:(f[275]>0)?276:(f[276]>0)?277:(f[277]>0)?278:(f[278]>0)?279:(f[279]>0)?280:(f[280]>0)?281:(f[281]>0)?282:(f[282]>0)?283:(f[283]>0)?284:(f[284]>0)?285:(f[285]>0)?286:(f[286]>0)?287:(f[287]>0)?288:(f[288]>0)?289:(f[289]>0)?290:(f[290]>0)?291:(f[291]>0)?292:(f[292]>0)?293:(f[293]>0)?294:(f[294]>0)?295:(f[295]>0)?296:(f[296]>0)?297:(f[297]>0)?298:(f[298]>0)?299:(f[299]>0)?300:(f[300]>0)?301:(f[301]>0)?302:(f[302]>0)?303:(f[303]>0)?304:(f[304]>0)?305:(f[305]>0)?306:(f[306]>0)?307:(f[307]>0)?308:(f[308]>0)?309:(f[309]>0)?310:(f[310]>0)?311:(f[311]>0)?312:(f[312]>0)?313:(f[313]>0)?314:(f[314]>0)?315:(f[315]>0)?316:(f[316]>0)?317:(f[317]>0)?318:(f[318]>0)?319:(f[319]>0)?320:(f[320]>0)?321:(f[321]>0)?322:(f[322]>0)?323:(f[323]>0)?324:(f[324]>0)?325:(f[325]>0)?326:(f[326]>0)?327:(f[327]>0)?328:(f[328]>0)?329:(f[329]>0)?330:(f[330]>0)?331:(f[331]>0)?332:(f[332]>0)?333:(f[333]>0)?334:(f[334]>0)?335:(f[335]>0)?336:(f[336]>0)?337:(f[337]>0)?338:(f[338]>0)?339:(f[339]>0)?340:(f[340]>0)?341:(f[341]>0)?342:(f[342]>0)?343:(f[343]>0)?344:(f[344]>0)?345:(f[345]>0)?346:(f[346]>0)?347:(f[347]>0)?348:(f[348]>0)?349:(f[349]>0)?350:(f[350]>0)?351:(f[351]>0)?352:(f[352]>0)?353:(f[353]>0)?354:(f[354]>0)?355:(f[355]>0)?356:(f[356]>0)?357:(f[357]>0)?358:(f[358]>0)?359:(f[359]>0)?360:(f[360]>0)?361:(f[361]>0)?362:(f[362]>0)?363:(f[363]>0)?364:(f[364]>0)?365:(f[365]>0)?366:(f[366]>0)?367:(f[367]>0)?368:(f[368]>0)?369:(f[369]>0)?370:(f[370]>0)?371:(f[371]>0)?372:(f[372]>0)?373:(f[373]>0)?374:(f[374]>0)?375:(f[375]>0)?376:(f[376]>0)?377:(f[377]>0)?378:(f[378]>0)?379:(f[379]>0)?380:(f[380]>0)?381:(f[381]>0)?382:(f[382]>0)?383:(f[383]>0)?384:(f[384]>0)?385:(f[385]>0)?386:(f[386]>0)?387:(f[387]>0)?388:(f[388]>0)?389:(f[389]>0)?390:(f[390]>0)?391:(f[391]>0)?392:(f[392]>0)?393:(f[393]>0)?394:(f[394]>0)?395:(f[395]>0)?396:(f[396]>0)?397:(f[397]>0)?398:(f[398]>0)?399:(f[399]>0)?400:(f[400]>0)?401:(f[401]>0)?402:(f[402]>0)?403:(f[403]>0)?404:(f[404]>0)?405:(f[405]>0)?406:(f[406]>0)?407:(f[407]>0)?408:(f[408]>0)?409:(f[409]>0)?410:(f[410]>0)?411:(f[411]>0)?412:(f[412]>0)?413:(f[413]>0)?414:(f[414]>0)?415:(f[415]>0)?416:(f[416]>0)?417:(f[417]>0)?418:(f[418]>0)?419:(f[419]>0)?420:(f[420]>0)?421:(f[421]>0)?422:(f[422]>0)?423:(f[423]>0)?424:(f[424]>0)?425:(f[425]>0)?426:(f[426]>0)?427:(f[427]>0)?428:(f[428]>0)?429:(f[429]>0)?430:(f[430]>0)?431:(f[431]>0)?432:(f[432]>0)?433:(f[433]>0)?434:(f[434]>0)?435:(f[435]>0)?436:(f[436]>0)?437:(f[437]>0)?438:(f[438]>0)?439:(f[439]>0)?440:(f[440]>0)?441:(f[441]>0)?442:(f[442]>0)?443:(f[443]>0)?444:(f[444]>0)?445:(f[445]>0)?446:(f[446]>0)?447:(f[447]>0)?448:(f[448]>0)?449:(f[449]>0)?450:(f[450]>0)?451:(f[451]>0)?452:(f[452]>0)?453:(f[453]>0)?454:(f[454]>0)?455:(f[455]>0)?456:(f[456]>0)?457:(f[457]>0)?458:(f[458]>0)?459:(f[459]>0)?460:(f[460]>0)?461:(f[461]>0)?462:(f[462]>0)?463:(f[463]>0)?464:(f[464]>0)?465:(f[465]>0)?466:(f[466]>0)?467:(f[467]>0)?468:(f[468]>0)?469:(f[469]>0)?470:(f[470]>0)?471:(f[471]>0)?472:(f[472]>0)?473:(f[473]>0)?474:(f[474]>0)?475:(f[475]>0)?476:(f[476]>0)?477:(f[477]>0)?478:(f[478]>0)?479:(f[479]>0)?480:(f[480]>0)?481:(f[481]>0)?482:(f[482]>0)?483:(f[483]>0)?484:(f[484]>0)?485:(f[485]>0)?486:(f[486]>0)?487:(f[487]>0)?488:(f[488]>0)?489:(f[489]>0)?490:(f[490]>0)?491:(f[491]>0)?492:(f[492]>0)?493:(f[493]>0)?494:(f[494]>0)?495:(f[495]>0)?496:(f[496]>0)?497:(f[497]>0)?498:(f[498]>0)?499:(f[499]>0)?500:(f[500]>0)?501:(f[501]>0)?502:(f[502]>0)?503:(f[503]>0)?504:(f[504]>0)?505:(f[505]>0)?506:(f[506]>0)?507:(f[507]>0)?508:(f[508]>0)?509:(f[509]>0)?510:(f[510]>0)?511:(f[511]>0)?512:(f[512]>0)?513:(f[513]>0)?514:(f[514]>0)?515:(f[515]>0)?516:(f[516]>0)?517:(f[517]>0)?518:(f[518]>0)?519:(f[519]>0)?520:(f[520]>0)?521:(f[521]>0)?522:(f[522]>0)?523:(f[523]>0)?524:(f[524]>0)?525:(f[525]>0)?526:(f[526]>0)?527:(f[527]>0)?528:(f[528]>0)?529:(f[529]>0)?530:(f[530]>0)?531:(f[531]>0)?532:(f[532]>0)?533:(f[533]>0)?534:(f[534]>0)?535:(f[535]>0)?536:(f[536]>0)?537:(f[537]>0)?538:(f[538]>0)?539:(f[539]>0)?540:(f[540]>0)?541:(f[541]>0)?542:(f[542]>0)?543:(f[543]>0)?544:(f[544]>0)?545:(f[545]>0)?546:(f[546]>0)?547:(f[547]>0)?548:(f[548]>0)?549:(f[549]>0)?550:(f[550]>0)?551:(f[551]>0)?552:(f[552]>0)?553:(f[553]>0)?554:(f[554]>0)?555:(f[555]>0)?556:(f[556]>0)?557:(f[557]>0)?558:(f[558]>0)?559:(f[559]>0)?560:(f[560]>0)?561:(f[561]>0)?562:(f[562]>0)?563:(f[563]>0)?564:(f[564]>0)?565:(f[565]>0)?566:(f[566]>0)?567:(f[567]>0)?568:(f[568]>0)?569:(f[569]>0)?570:(f[570]>0)?571:(f[571]>0)?572:(f[572]>0)?573:(f[573]>0)?574:(f[574]>0)?575:(f[575]>0)?576:(f[576]>0)?577:(f[577]>0)?578:(f[578]>0)?579:(f[579]>0)?580:(f[580]>0)?581:(f[581]>0)?582:(f[582]>0)?583:(f[583]>0)?584:(f[584]>0)?585:(f[585]>0)?586:(f[586]>0)?587:(f[587]>0)?588:(f[588]>0)?589:(f[589]>0)?590:(f[590]>0)?591:(f[591]>0)?592:(f[592]>0)?593:(f[593]>0)?594:(f[594]>0)?595:(f[595]>0)?596:(f[596]>0)?597:(f[597]>0)?598:(f[598]>0)?599:(f[599]>0)?600:(f[600]>0)?601:(f[601]>0)?602:(f[602]>0)?603:(f[603]>0)?604:(f[604]>0)?605:(f[605]>0)?606:(f[606]>0)?607:(f[607]>0)?608:(f[608]>0)?609:(f[609]>0)?610:(f[610]>0)?611:(f[611]>0)?612:(f[612]>0)?613:(f[613]>0)?614:(f[614]>0)?615:(f[615]>0)?616:(f[616]>0)?617:(f[617]>0)?618:(f[618]>0)?619:(f[619]>0)?620:(f[620]>0)?621:(f[621]>0)?622:(f[622]>0)?623:(f[623]>0)?624:(f[624]>0)?625:(f[625]>0)?626:(f[626]>0)?627:(f[627]>0)?628:(f[628]>0)?629:(f[629]>0)?630:(f[630]>0)?631:(f[631]>0)?632:(f[632]>0)?633:(f[633]>0)?634:(f[634]>0)?635:(f[635]>0)?636:(f[636]>0)?637:(f[637]>0)?638:(f[638]>0)?639:(f[639]>0)?640:(f[640]>0)?641:(f[641]>0)?642:(f[642]>0)?643:(f[643]>0)?644:(f[644]>0)?645:(f[645]>0)?646:(f[646]>0)?647:(f[647]>0)?648:(f[648]>0)?649:(f[649]>0)?650:(f[650]>0)?651:(f[651]>0)?652:(f[652]>0)?653:(f[653]>0)?654:(f[654]>0)?655:(f[655]>0)?656:(f[656]>0)?657:(f[657]>0)?658:(f[658]>0)?659:(f[659]>0)?660:(f[660]>0)?661:(f[661]>0)?662:(f[662]>0)?663:(f[663]>0)?664:(f[664]>0)?665:(f[665]>0)?666:(f[666]>0)?667:(f[667]>0)?668:(f[668]>0)?669:(f[669]>0)?670:(f[670]>0)?671:(f[671]>0)?672:(f[672]>0)?673:(f[673]>0)?674:(f[674]>0)?675:(f[675]>0)?676:(f[676]>0)?677:(f[677]>0)?678:(f[678]>0)?679:(f[679]>0)?680:(f[680]>0)?681:(f[681]>0)?682:(f[682]>0)?683:(f[683]>0)?684:(f[684]>0)?685:(f[685]>0)?686:(f[686]>0)?687:(f[687]>0)?688:(f[688]>0)?689:(f[689]>0)?690:(f[690]>0)?691:(f[691]>0)?692:(f[692]>0)?693:(f[693]>0)?694:(f[694]>0)?695:(f[695]>0)?696:(f[696]>0)?697:(f[697]>0)?698:(f[698]>0)?699:(f[699]>0)?700:(f[700]>0)?701:(f[701]>0)?702:(f[702]>0)?703:(f[703]>0)?704:(f[704]>0)?705:(f[705]>0)?706:(f[706]>0)?707:(f[707]>0)?708:(f[708]>0)?709:(f[709]>0)?710:(f[710]>0)?711:(f[711]>0)?712:(f[712]>0)?713:(f[713]>0)?714:(f[714]>0)?715:(f[715]>0)?716:(f[716]>0)?717:(f[717]>0)?718:(f[718]>0)?719:(f[719]>0)?720:(f[720]>0)?721:(f[721]>0)?722:(f[722]>0)?723:(f[723]>0)?724:(f[724]>0)?725:(f[725]>0)?726:(f[726]>0)?727:(f[727]>0)?728:(f[728]>0)?729:(f[729]>0)?730:(f[730]>0)?731:(f[731]>0)?732:0;
        case(tf)
                1: begin
                        tc = f[0];
                        p[88] = p[88] - tc;
                        p[85] = p[85] + tc;
                end
                2: begin
                        tc = f[1];
                        p[112] = p[112] - tc;
                        p[109] = p[109] + tc;
                end
                3: begin
                        tc = f[2];
                        p[136] = p[136] - tc;
                        p[133] = p[133] + tc;
                end
                4: begin
                        tc = f[3];
                        p[160] = p[160] - tc;
                        p[157] = p[157] + tc;
                end
                5: begin
                        tc = f[4];
                        p[184] = p[184] - tc;
                        p[181] = p[181] + tc;
                end
                6: begin
                        tc = f[5];
                        p[208] = p[208] - tc;
                        p[205] = p[205] + tc;
                end
                7: begin
                        tc = f[6];
                        p[232] = p[232] - tc;
                        p[229] = p[229] + tc;
                end
                8: begin
                        tc = f[7];
                        p[256] = p[256] - tc;
                        p[253] = p[253] + tc;
                end
                9: begin
                        tc = f[8];
                        p[280] = p[280] - tc;
                        p[277] = p[277] + tc;
                end
                10: begin
                        tc = f[9];
                        p[304] = p[304] - tc;
                        p[301] = p[301] + tc;
                end
                11: begin
                        tc = f[10];
                        p[328] = p[328] - tc;
                        p[325] = p[325] + tc;
                end
                12: begin
                        tc = f[11];
                        p[347] = p[347] - tc;
                        p[349] = p[349] + tc;
                end
                13: begin
                        tc = f[12];
                        p[366] = p[366] - tc;
                        p[363] = p[363] + tc;
                end
                14: begin
                        tc = f[13];
                        p[390] = p[390] - tc;
                        p[387] = p[387] + tc;
                end
                15: begin
                        tc = f[14];
                        p[414] = p[414] - tc;
                        p[411] = p[411] + tc;
                end
                16: begin
                        tc = f[15];
                        p[438] = p[438] - tc;
                        p[435] = p[435] + tc;
                end
                17: begin
                        tc = f[16];
                        p[457] = p[457] - tc;
                        p[459] = p[459] + tc;
                end
                18: begin
                        tc = f[17];
                        p[476] = p[476] - tc;
                        p[473] = p[473] + tc;
                end
                19: begin
                        tc = f[18];
                        p[500] = p[500] - tc;
                        p[497] = p[497] + tc;
                end
                20: begin
                        tc = f[19];
                        p[524] = p[524] - tc;
                        p[521] = p[521] + tc;
                end
                21: begin
                        tc = f[20];
                        p[543] = p[543] - tc;
                        p[545] = p[545] + tc;
                end
                22: begin
                        tc = f[21];
                        p[562] = p[562] - tc;
                        p[559] = p[559] + tc;
                end
                23: begin
                        tc = f[22];
                        p[586] = p[586] - tc;
                        p[583] = p[583] + tc;
                end
                24: begin
                        tc = f[23];
                        p[605] = p[605] - tc;
                        p[607] = p[607] + tc;
                end
                25: begin
                        tc = f[24];
                        p[624] = p[624] - tc;
                        p[621] = p[621] + tc;
                end
                26: begin
                        tc = f[25];
                        p[643] = p[643] - tc;
                        p[645] = p[645] + tc;
                end
                27: begin
                        tc = f[26];
                        p[657] = p[657] - tc;
                        p[659] = p[659] + tc;
                end
                28: begin
                        tc = f[27];
                        p[89] = p[89] - tc;
                        p[85] = p[85] + tc;
                end
                29: begin
                        tc = f[28];
                        p[83] = p[83] - tc;
                end
                30: begin
                        tc = f[29];
                        p[87] = p[87] - tc;
                        p[89] = p[89] + tc;
                end
                31: begin
                        tc = f[30];
                        p[84] = p[84] - tc*2;
                        p[90] = p[90] + tc;
                end
                32: begin
                        tc = f[31];
                        p[91] = p[91] - tc;
                        p[88] = p[88] + tc;
                end
                33: begin
                        tc = f[32];
                        p[84] = p[84] - tc;
                        p[93] = p[93] - tc;
                        p[92] = p[92] + tc;
                end
                34: begin
                        tc = f[33];
                        p[94] = p[94] - tc;
                        p[91] = p[91] + tc;
                end
                35: begin
                        tc = f[34];
                        p[83] = p[83] - tc;
                        p[86] = p[86] + tc;
                        p[95] = p[95] + tc;
                end
                36: begin
                        tc = f[35];
                        p[83] = p[83] - tc;
                        p[95] = p[95] + tc;
                end
                37: begin
                        tc = f[36];
                        p[96] = p[96] - tc;
                        p[94] = p[94] + tc;
                end
                38: begin
                        tc = f[37];
                        p[90] = p[90] - tc;
                        p[84] = p[84] + tc;
                end
                39: begin
                        tc = f[38];
                        p[97] = p[97] - tc;
                        p[96] = p[96] + tc;
                end
                40: begin
                        tc = f[39];
                        p[95] = p[95] - tc;
                        p[83] = p[83] + tc*2;
                end
                41: begin
                        tc = f[40];
                        p[85] = p[85] - tc;
                        p[92] = p[92] - tc;
                        p[93] = p[93] + tc;
                        p[97] = p[97] + tc;
                end
                42: begin
                        tc = f[41];
                        p[85] = p[85] - tc;
                        p[97] = p[97] + tc;
                end
                43: begin
                        tc = f[42];
                        p[28] = p[28] - tc;
                        p[83] = p[83] + tc;
                        p[98] = p[98] + tc;
                end
                44: begin
                        tc = f[43];
                        p[98] = p[98] - tc;
                        p[28] = p[28] + tc;
                end
                45: begin
                        tc = f[44];
                        p[100] = p[100] - tc;
                        p[99] = p[99] + tc;
                end
                46: begin
                        tc = f[45];
                        p[101] = p[101] - tc;
                        p[100] = p[100] + tc;
                end
                47: begin
                        tc = f[46];
                        p[29] = p[29] - tc;
                        p[84] = p[84] + tc;
                        p[102] = p[102] + tc;
                end
                48: begin
                        tc = f[47];
                        p[102] = p[102] - tc;
                        p[29] = p[29] + tc;
                end
                49: begin
                        tc = f[48];
                        p[104] = p[104] - tc;
                        p[103] = p[103] + tc;
                end
                50: begin
                        tc = f[49];
                        p[105] = p[105] - tc;
                        p[104] = p[104] + tc;
                end
                51: begin
                        tc = f[50];
                        p[99] = p[99] - tc;
                        p[103] = p[103] - tc;
                        p[0] = p[0] + tc;
                end
                52: begin
                        tc = f[51];
                        p[85] = p[85] - tc;
                        p[101] = p[101] + tc;
                        p[105] = p[105] + tc;
                end
                53: begin
                        tc = f[52];
                        p[86] = p[86] - tc;
                        p[30] = p[30] + tc;
                end
                54: begin
                        tc = f[53];
                        p[30] = p[30] - tc;
                end
                55: begin
                        tc = f[54];
                        p[106] = p[106] - tc;
                        p[87] = p[87] + tc;
                end
                56: begin
                        tc = f[55];
                        p[1] = p[1] - tc;
                        p[106] = p[106] + tc;
                end
                57: begin
                        tc = f[56];
                        p[113] = p[113] - tc;
                        p[109] = p[109] + tc;
                end
                58: begin
                        tc = f[57];
                        p[107] = p[107] - tc;
                end
                59: begin
                        tc = f[58];
                        p[111] = p[111] - tc;
                        p[113] = p[113] + tc;
                end
                60: begin
                        tc = f[59];
                        p[108] = p[108] - tc*2;
                        p[114] = p[114] + tc;
                end
                61: begin
                        tc = f[60];
                        p[115] = p[115] - tc;
                        p[112] = p[112] + tc;
                end
                62: begin
                        tc = f[61];
                        p[108] = p[108] - tc;
                        p[117] = p[117] - tc;
                        p[116] = p[116] + tc;
                end
                63: begin
                        tc = f[62];
                        p[118] = p[118] - tc;
                        p[115] = p[115] + tc;
                end
                64: begin
                        tc = f[63];
                        p[107] = p[107] - tc;
                        p[110] = p[110] + tc;
                        p[119] = p[119] + tc;
                end
                65: begin
                        tc = f[64];
                        p[107] = p[107] - tc;
                        p[119] = p[119] + tc;
                end
                66: begin
                        tc = f[65];
                        p[120] = p[120] - tc;
                        p[118] = p[118] + tc;
                end
                67: begin
                        tc = f[66];
                        p[114] = p[114] - tc;
                        p[108] = p[108] + tc;
                end
                68: begin
                        tc = f[67];
                        p[121] = p[121] - tc;
                        p[120] = p[120] + tc;
                end
                69: begin
                        tc = f[68];
                        p[119] = p[119] - tc;
                        p[107] = p[107] + tc*2;
                end
                70: begin
                        tc = f[69];
                        p[109] = p[109] - tc;
                        p[116] = p[116] - tc;
                        p[117] = p[117] + tc;
                        p[121] = p[121] + tc;
                end
                71: begin
                        tc = f[70];
                        p[109] = p[109] - tc;
                        p[121] = p[121] + tc;
                end
                72: begin
                        tc = f[71];
                        p[30] = p[30] - tc;
                        p[107] = p[107] + tc;
                        p[122] = p[122] + tc;
                end
                73: begin
                        tc = f[72];
                        p[122] = p[122] - tc;
                        p[30] = p[30] + tc;
                end
                74: begin
                        tc = f[73];
                        p[124] = p[124] - tc;
                        p[123] = p[123] + tc;
                end
                75: begin
                        tc = f[74];
                        p[125] = p[125] - tc;
                        p[124] = p[124] + tc;
                end
                76: begin
                        tc = f[75];
                        p[31] = p[31] - tc;
                        p[108] = p[108] + tc;
                        p[126] = p[126] + tc;
                end
                77: begin
                        tc = f[76];
                        p[126] = p[126] - tc;
                        p[31] = p[31] + tc;
                end
                78: begin
                        tc = f[77];
                        p[128] = p[128] - tc;
                        p[127] = p[127] + tc;
                end
                79: begin
                        tc = f[78];
                        p[129] = p[129] - tc;
                        p[128] = p[128] + tc;
                end
                80: begin
                        tc = f[79];
                        p[123] = p[123] - tc;
                        p[127] = p[127] - tc;
                        p[1] = p[1] + tc;
                end
                81: begin
                        tc = f[80];
                        p[109] = p[109] - tc;
                        p[125] = p[125] + tc;
                        p[129] = p[129] + tc;
                end
                82: begin
                        tc = f[81];
                        p[110] = p[110] - tc;
                        p[32] = p[32] + tc;
                end
                83: begin
                        tc = f[82];
                        p[32] = p[32] - tc;
                end
                84: begin
                        tc = f[83];
                        p[130] = p[130] - tc;
                        p[111] = p[111] + tc;
                end
                85: begin
                        tc = f[84];
                        p[2] = p[2] - tc;
                        p[130] = p[130] + tc;
                end
                86: begin
                        tc = f[85];
                        p[137] = p[137] - tc;
                        p[133] = p[133] + tc;
                end
                87: begin
                        tc = f[86];
                        p[131] = p[131] - tc;
                end
                88: begin
                        tc = f[87];
                        p[135] = p[135] - tc;
                        p[137] = p[137] + tc;
                end
                89: begin
                        tc = f[88];
                        p[132] = p[132] - tc*2;
                        p[138] = p[138] + tc;
                end
                90: begin
                        tc = f[89];
                        p[139] = p[139] - tc;
                        p[136] = p[136] + tc;
                end
                91: begin
                        tc = f[90];
                        p[132] = p[132] - tc;
                        p[141] = p[141] - tc;
                        p[140] = p[140] + tc;
                end
                92: begin
                        tc = f[91];
                        p[142] = p[142] - tc;
                        p[139] = p[139] + tc;
                end
                93: begin
                        tc = f[92];
                        p[131] = p[131] - tc;
                        p[134] = p[134] + tc;
                        p[143] = p[143] + tc;
                end
                94: begin
                        tc = f[93];
                        p[131] = p[131] - tc;
                        p[143] = p[143] + tc;
                end
                95: begin
                        tc = f[94];
                        p[144] = p[144] - tc;
                        p[142] = p[142] + tc;
                end
                96: begin
                        tc = f[95];
                        p[138] = p[138] - tc;
                        p[132] = p[132] + tc;
                end
                97: begin
                        tc = f[96];
                        p[145] = p[145] - tc;
                        p[144] = p[144] + tc;
                end
                98: begin
                        tc = f[97];
                        p[143] = p[143] - tc;
                        p[131] = p[131] + tc*2;
                end
                99: begin
                        tc = f[98];
                        p[133] = p[133] - tc;
                        p[140] = p[140] - tc;
                        p[141] = p[141] + tc;
                        p[145] = p[145] + tc;
                end
                100: begin
                        tc = f[99];
                        p[133] = p[133] - tc;
                        p[145] = p[145] + tc;
                end
                101: begin
                        tc = f[100];
                        p[32] = p[32] - tc;
                        p[131] = p[131] + tc;
                        p[146] = p[146] + tc;
                end
                102: begin
                        tc = f[101];
                        p[146] = p[146] - tc;
                        p[32] = p[32] + tc;
                end
                103: begin
                        tc = f[102];
                        p[148] = p[148] - tc;
                        p[147] = p[147] + tc;
                end
                104: begin
                        tc = f[103];
                        p[149] = p[149] - tc;
                        p[148] = p[148] + tc;
                end
                105: begin
                        tc = f[104];
                        p[33] = p[33] - tc;
                        p[132] = p[132] + tc;
                        p[150] = p[150] + tc;
                end
                106: begin
                        tc = f[105];
                        p[150] = p[150] - tc;
                        p[33] = p[33] + tc;
                end
                107: begin
                        tc = f[106];
                        p[152] = p[152] - tc;
                        p[151] = p[151] + tc;
                end
                108: begin
                        tc = f[107];
                        p[153] = p[153] - tc;
                        p[152] = p[152] + tc;
                end
                109: begin
                        tc = f[108];
                        p[147] = p[147] - tc;
                        p[151] = p[151] - tc;
                        p[2] = p[2] + tc;
                end
                110: begin
                        tc = f[109];
                        p[133] = p[133] - tc;
                        p[149] = p[149] + tc;
                        p[153] = p[153] + tc;
                end
                111: begin
                        tc = f[110];
                        p[134] = p[134] - tc;
                        p[34] = p[34] + tc;
                end
                112: begin
                        tc = f[111];
                        p[34] = p[34] - tc;
                end
                113: begin
                        tc = f[112];
                        p[154] = p[154] - tc;
                        p[135] = p[135] + tc;
                end
                114: begin
                        tc = f[113];
                        p[3] = p[3] - tc;
                        p[154] = p[154] + tc;
                end
                115: begin
                        tc = f[114];
                        p[161] = p[161] - tc;
                        p[157] = p[157] + tc;
                end
                116: begin
                        tc = f[115];
                        p[155] = p[155] - tc;
                end
                117: begin
                        tc = f[116];
                        p[159] = p[159] - tc;
                        p[161] = p[161] + tc;
                end
                118: begin
                        tc = f[117];
                        p[156] = p[156] - tc*2;
                        p[162] = p[162] + tc;
                end
                119: begin
                        tc = f[118];
                        p[163] = p[163] - tc;
                        p[160] = p[160] + tc;
                end
                120: begin
                        tc = f[119];
                        p[156] = p[156] - tc;
                        p[165] = p[165] - tc;
                        p[164] = p[164] + tc;
                end
                121: begin
                        tc = f[120];
                        p[166] = p[166] - tc;
                        p[163] = p[163] + tc;
                end
                122: begin
                        tc = f[121];
                        p[155] = p[155] - tc;
                        p[158] = p[158] + tc;
                        p[167] = p[167] + tc;
                end
                123: begin
                        tc = f[122];
                        p[155] = p[155] - tc;
                        p[167] = p[167] + tc;
                end
                124: begin
                        tc = f[123];
                        p[168] = p[168] - tc;
                        p[166] = p[166] + tc;
                end
                125: begin
                        tc = f[124];
                        p[162] = p[162] - tc;
                        p[156] = p[156] + tc;
                end
                126: begin
                        tc = f[125];
                        p[169] = p[169] - tc;
                        p[168] = p[168] + tc;
                end
                127: begin
                        tc = f[126];
                        p[167] = p[167] - tc;
                        p[155] = p[155] + tc*2;
                end
                128: begin
                        tc = f[127];
                        p[157] = p[157] - tc;
                        p[164] = p[164] - tc;
                        p[165] = p[165] + tc;
                        p[169] = p[169] + tc;
                end
                129: begin
                        tc = f[128];
                        p[157] = p[157] - tc;
                        p[169] = p[169] + tc;
                end
                130: begin
                        tc = f[129];
                        p[34] = p[34] - tc;
                        p[155] = p[155] + tc;
                        p[170] = p[170] + tc;
                end
                131: begin
                        tc = f[130];
                        p[170] = p[170] - tc;
                        p[34] = p[34] + tc;
                end
                132: begin
                        tc = f[131];
                        p[172] = p[172] - tc;
                        p[171] = p[171] + tc;
                end
                133: begin
                        tc = f[132];
                        p[173] = p[173] - tc;
                        p[172] = p[172] + tc;
                end
                134: begin
                        tc = f[133];
                        p[35] = p[35] - tc;
                        p[156] = p[156] + tc;
                        p[174] = p[174] + tc;
                end
                135: begin
                        tc = f[134];
                        p[174] = p[174] - tc;
                        p[35] = p[35] + tc;
                end
                136: begin
                        tc = f[135];
                        p[176] = p[176] - tc;
                        p[175] = p[175] + tc;
                end
                137: begin
                        tc = f[136];
                        p[177] = p[177] - tc;
                        p[176] = p[176] + tc;
                end
                138: begin
                        tc = f[137];
                        p[171] = p[171] - tc;
                        p[175] = p[175] - tc;
                        p[3] = p[3] + tc;
                end
                139: begin
                        tc = f[138];
                        p[157] = p[157] - tc;
                        p[173] = p[173] + tc;
                        p[177] = p[177] + tc;
                end
                140: begin
                        tc = f[139];
                        p[158] = p[158] - tc;
                        p[36] = p[36] + tc;
                end
                141: begin
                        tc = f[140];
                        p[36] = p[36] - tc;
                end
                142: begin
                        tc = f[141];
                        p[178] = p[178] - tc;
                        p[159] = p[159] + tc;
                end
                143: begin
                        tc = f[142];
                        p[4] = p[4] - tc;
                        p[178] = p[178] + tc;
                end
                144: begin
                        tc = f[143];
                        p[185] = p[185] - tc;
                        p[181] = p[181] + tc;
                end
                145: begin
                        tc = f[144];
                        p[179] = p[179] - tc;
                end
                146: begin
                        tc = f[145];
                        p[183] = p[183] - tc;
                        p[185] = p[185] + tc;
                end
                147: begin
                        tc = f[146];
                        p[180] = p[180] - tc*2;
                        p[186] = p[186] + tc;
                end
                148: begin
                        tc = f[147];
                        p[187] = p[187] - tc;
                        p[184] = p[184] + tc;
                end
                149: begin
                        tc = f[148];
                        p[180] = p[180] - tc;
                        p[189] = p[189] - tc;
                        p[188] = p[188] + tc;
                end
                150: begin
                        tc = f[149];
                        p[190] = p[190] - tc;
                        p[187] = p[187] + tc;
                end
                151: begin
                        tc = f[150];
                        p[179] = p[179] - tc;
                        p[182] = p[182] + tc;
                        p[191] = p[191] + tc;
                end
                152: begin
                        tc = f[151];
                        p[179] = p[179] - tc;
                        p[191] = p[191] + tc;
                end
                153: begin
                        tc = f[152];
                        p[192] = p[192] - tc;
                        p[190] = p[190] + tc;
                end
                154: begin
                        tc = f[153];
                        p[186] = p[186] - tc;
                        p[180] = p[180] + tc;
                end
                155: begin
                        tc = f[154];
                        p[193] = p[193] - tc;
                        p[192] = p[192] + tc;
                end
                156: begin
                        tc = f[155];
                        p[191] = p[191] - tc;
                        p[179] = p[179] + tc*2;
                end
                157: begin
                        tc = f[156];
                        p[181] = p[181] - tc;
                        p[188] = p[188] - tc;
                        p[189] = p[189] + tc;
                        p[193] = p[193] + tc;
                end
                158: begin
                        tc = f[157];
                        p[181] = p[181] - tc;
                        p[193] = p[193] + tc;
                end
                159: begin
                        tc = f[158];
                        p[36] = p[36] - tc;
                        p[179] = p[179] + tc;
                        p[194] = p[194] + tc;
                end
                160: begin
                        tc = f[159];
                        p[194] = p[194] - tc;
                        p[36] = p[36] + tc;
                end
                161: begin
                        tc = f[160];
                        p[196] = p[196] - tc;
                        p[195] = p[195] + tc;
                end
                162: begin
                        tc = f[161];
                        p[197] = p[197] - tc;
                        p[196] = p[196] + tc;
                end
                163: begin
                        tc = f[162];
                        p[37] = p[37] - tc;
                        p[180] = p[180] + tc;
                        p[198] = p[198] + tc;
                end
                164: begin
                        tc = f[163];
                        p[198] = p[198] - tc;
                        p[37] = p[37] + tc;
                end
                165: begin
                        tc = f[164];
                        p[200] = p[200] - tc;
                        p[199] = p[199] + tc;
                end
                166: begin
                        tc = f[165];
                        p[201] = p[201] - tc;
                        p[200] = p[200] + tc;
                end
                167: begin
                        tc = f[166];
                        p[195] = p[195] - tc;
                        p[199] = p[199] - tc;
                        p[4] = p[4] + tc;
                end
                168: begin
                        tc = f[167];
                        p[181] = p[181] - tc;
                        p[197] = p[197] + tc;
                        p[201] = p[201] + tc;
                end
                169: begin
                        tc = f[168];
                        p[182] = p[182] - tc;
                        p[38] = p[38] + tc;
                end
                170: begin
                        tc = f[169];
                        p[38] = p[38] - tc;
                end
                171: begin
                        tc = f[170];
                        p[202] = p[202] - tc;
                        p[183] = p[183] + tc;
                end
                172: begin
                        tc = f[171];
                        p[5] = p[5] - tc;
                        p[202] = p[202] + tc;
                end
                173: begin
                        tc = f[172];
                        p[209] = p[209] - tc;
                        p[205] = p[205] + tc;
                end
                174: begin
                        tc = f[173];
                        p[203] = p[203] - tc;
                end
                175: begin
                        tc = f[174];
                        p[207] = p[207] - tc;
                        p[209] = p[209] + tc;
                end
                176: begin
                        tc = f[175];
                        p[204] = p[204] - tc*2;
                        p[210] = p[210] + tc;
                end
                177: begin
                        tc = f[176];
                        p[211] = p[211] - tc;
                        p[208] = p[208] + tc;
                end
                178: begin
                        tc = f[177];
                        p[204] = p[204] - tc;
                        p[213] = p[213] - tc;
                        p[212] = p[212] + tc;
                end
                179: begin
                        tc = f[178];
                        p[214] = p[214] - tc;
                        p[211] = p[211] + tc;
                end
                180: begin
                        tc = f[179];
                        p[203] = p[203] - tc;
                        p[206] = p[206] + tc;
                        p[215] = p[215] + tc;
                end
                181: begin
                        tc = f[180];
                        p[203] = p[203] - tc;
                        p[215] = p[215] + tc;
                end
                182: begin
                        tc = f[181];
                        p[216] = p[216] - tc;
                        p[214] = p[214] + tc;
                end
                183: begin
                        tc = f[182];
                        p[210] = p[210] - tc;
                        p[204] = p[204] + tc;
                end
                184: begin
                        tc = f[183];
                        p[217] = p[217] - tc;
                        p[216] = p[216] + tc;
                end
                185: begin
                        tc = f[184];
                        p[215] = p[215] - tc;
                        p[203] = p[203] + tc*2;
                end
                186: begin
                        tc = f[185];
                        p[205] = p[205] - tc;
                        p[212] = p[212] - tc;
                        p[213] = p[213] + tc;
                        p[217] = p[217] + tc;
                end
                187: begin
                        tc = f[186];
                        p[205] = p[205] - tc;
                        p[217] = p[217] + tc;
                end
                188: begin
                        tc = f[187];
                        p[38] = p[38] - tc;
                        p[203] = p[203] + tc;
                        p[218] = p[218] + tc;
                end
                189: begin
                        tc = f[188];
                        p[218] = p[218] - tc;
                        p[38] = p[38] + tc;
                end
                190: begin
                        tc = f[189];
                        p[220] = p[220] - tc;
                        p[219] = p[219] + tc;
                end
                191: begin
                        tc = f[190];
                        p[221] = p[221] - tc;
                        p[220] = p[220] + tc;
                end
                192: begin
                        tc = f[191];
                        p[39] = p[39] - tc;
                        p[204] = p[204] + tc;
                        p[222] = p[222] + tc;
                end
                193: begin
                        tc = f[192];
                        p[222] = p[222] - tc;
                        p[39] = p[39] + tc;
                end
                194: begin
                        tc = f[193];
                        p[224] = p[224] - tc;
                        p[223] = p[223] + tc;
                end
                195: begin
                        tc = f[194];
                        p[225] = p[225] - tc;
                        p[224] = p[224] + tc;
                end
                196: begin
                        tc = f[195];
                        p[219] = p[219] - tc;
                        p[223] = p[223] - tc;
                        p[5] = p[5] + tc;
                end
                197: begin
                        tc = f[196];
                        p[205] = p[205] - tc;
                        p[221] = p[221] + tc;
                        p[225] = p[225] + tc;
                end
                198: begin
                        tc = f[197];
                        p[206] = p[206] - tc;
                        p[40] = p[40] + tc;
                end
                199: begin
                        tc = f[198];
                        p[40] = p[40] - tc;
                end
                200: begin
                        tc = f[199];
                        p[226] = p[226] - tc;
                        p[207] = p[207] + tc;
                end
                201: begin
                        tc = f[200];
                        p[6] = p[6] - tc;
                        p[226] = p[226] + tc;
                end
                202: begin
                        tc = f[201];
                        p[233] = p[233] - tc;
                        p[229] = p[229] + tc;
                end
                203: begin
                        tc = f[202];
                        p[227] = p[227] - tc;
                end
                204: begin
                        tc = f[203];
                        p[231] = p[231] - tc;
                        p[233] = p[233] + tc;
                end
                205: begin
                        tc = f[204];
                        p[228] = p[228] - tc*2;
                        p[234] = p[234] + tc;
                end
                206: begin
                        tc = f[205];
                        p[235] = p[235] - tc;
                        p[232] = p[232] + tc;
                end
                207: begin
                        tc = f[206];
                        p[228] = p[228] - tc;
                        p[237] = p[237] - tc;
                        p[236] = p[236] + tc;
                end
                208: begin
                        tc = f[207];
                        p[238] = p[238] - tc;
                        p[235] = p[235] + tc;
                end
                209: begin
                        tc = f[208];
                        p[227] = p[227] - tc;
                        p[230] = p[230] + tc;
                        p[239] = p[239] + tc;
                end
                210: begin
                        tc = f[209];
                        p[227] = p[227] - tc;
                        p[239] = p[239] + tc;
                end
                211: begin
                        tc = f[210];
                        p[240] = p[240] - tc;
                        p[238] = p[238] + tc;
                end
                212: begin
                        tc = f[211];
                        p[234] = p[234] - tc;
                        p[228] = p[228] + tc;
                end
                213: begin
                        tc = f[212];
                        p[241] = p[241] - tc;
                        p[240] = p[240] + tc;
                end
                214: begin
                        tc = f[213];
                        p[239] = p[239] - tc;
                        p[227] = p[227] + tc*2;
                end
                215: begin
                        tc = f[214];
                        p[229] = p[229] - tc;
                        p[236] = p[236] - tc;
                        p[237] = p[237] + tc;
                        p[241] = p[241] + tc;
                end
                216: begin
                        tc = f[215];
                        p[229] = p[229] - tc;
                        p[241] = p[241] + tc;
                end
                217: begin
                        tc = f[216];
                        p[41] = p[41] - tc;
                        p[227] = p[227] + tc;
                        p[242] = p[242] + tc;
                end
                218: begin
                        tc = f[217];
                        p[242] = p[242] - tc;
                        p[41] = p[41] + tc;
                end
                219: begin
                        tc = f[218];
                        p[244] = p[244] - tc;
                        p[243] = p[243] + tc;
                end
                220: begin
                        tc = f[219];
                        p[245] = p[245] - tc;
                        p[244] = p[244] + tc;
                end
                221: begin
                        tc = f[220];
                        p[42] = p[42] - tc;
                        p[228] = p[228] + tc;
                        p[246] = p[246] + tc;
                end
                222: begin
                        tc = f[221];
                        p[246] = p[246] - tc;
                        p[42] = p[42] + tc;
                end
                223: begin
                        tc = f[222];
                        p[248] = p[248] - tc;
                        p[247] = p[247] + tc;
                end
                224: begin
                        tc = f[223];
                        p[249] = p[249] - tc;
                        p[248] = p[248] + tc;
                end
                225: begin
                        tc = f[224];
                        p[243] = p[243] - tc;
                        p[247] = p[247] - tc;
                        p[6] = p[6] + tc;
                end
                226: begin
                        tc = f[225];
                        p[229] = p[229] - tc;
                        p[245] = p[245] + tc;
                        p[249] = p[249] + tc;
                end
                227: begin
                        tc = f[226];
                        p[230] = p[230] - tc;
                        p[43] = p[43] + tc;
                end
                228: begin
                        tc = f[227];
                        p[43] = p[43] - tc;
                end
                229: begin
                        tc = f[228];
                        p[250] = p[250] - tc;
                        p[231] = p[231] + tc;
                end
                230: begin
                        tc = f[229];
                        p[7] = p[7] - tc;
                        p[250] = p[250] + tc;
                end
                231: begin
                        tc = f[230];
                        p[257] = p[257] - tc;
                        p[253] = p[253] + tc;
                end
                232: begin
                        tc = f[231];
                        p[251] = p[251] - tc;
                end
                233: begin
                        tc = f[232];
                        p[255] = p[255] - tc;
                        p[257] = p[257] + tc;
                end
                234: begin
                        tc = f[233];
                        p[252] = p[252] - tc*2;
                        p[258] = p[258] + tc;
                end
                235: begin
                        tc = f[234];
                        p[259] = p[259] - tc;
                        p[256] = p[256] + tc;
                end
                236: begin
                        tc = f[235];
                        p[252] = p[252] - tc;
                        p[261] = p[261] - tc;
                        p[260] = p[260] + tc;
                end
                237: begin
                        tc = f[236];
                        p[262] = p[262] - tc;
                        p[259] = p[259] + tc;
                end
                238: begin
                        tc = f[237];
                        p[251] = p[251] - tc;
                        p[254] = p[254] + tc;
                        p[263] = p[263] + tc;
                end
                239: begin
                        tc = f[238];
                        p[251] = p[251] - tc;
                        p[263] = p[263] + tc;
                end
                240: begin
                        tc = f[239];
                        p[264] = p[264] - tc;
                        p[262] = p[262] + tc;
                end
                241: begin
                        tc = f[240];
                        p[258] = p[258] - tc;
                        p[252] = p[252] + tc;
                end
                242: begin
                        tc = f[241];
                        p[265] = p[265] - tc;
                        p[264] = p[264] + tc;
                end
                243: begin
                        tc = f[242];
                        p[263] = p[263] - tc;
                        p[251] = p[251] + tc*2;
                end
                244: begin
                        tc = f[243];
                        p[253] = p[253] - tc;
                        p[260] = p[260] - tc;
                        p[261] = p[261] + tc;
                        p[265] = p[265] + tc;
                end
                245: begin
                        tc = f[244];
                        p[253] = p[253] - tc;
                        p[265] = p[265] + tc;
                end
                246: begin
                        tc = f[245];
                        p[43] = p[43] - tc;
                        p[251] = p[251] + tc;
                        p[266] = p[266] + tc;
                end
                247: begin
                        tc = f[246];
                        p[266] = p[266] - tc;
                        p[43] = p[43] + tc;
                end
                248: begin
                        tc = f[247];
                        p[268] = p[268] - tc;
                        p[267] = p[267] + tc;
                end
                249: begin
                        tc = f[248];
                        p[269] = p[269] - tc;
                        p[268] = p[268] + tc;
                end
                250: begin
                        tc = f[249];
                        p[44] = p[44] - tc;
                        p[252] = p[252] + tc;
                        p[270] = p[270] + tc;
                end
                251: begin
                        tc = f[250];
                        p[270] = p[270] - tc;
                        p[44] = p[44] + tc;
                end
                252: begin
                        tc = f[251];
                        p[272] = p[272] - tc;
                        p[271] = p[271] + tc;
                end
                253: begin
                        tc = f[252];
                        p[273] = p[273] - tc;
                        p[272] = p[272] + tc;
                end
                254: begin
                        tc = f[253];
                        p[267] = p[267] - tc;
                        p[271] = p[271] - tc;
                        p[7] = p[7] + tc;
                end
                255: begin
                        tc = f[254];
                        p[253] = p[253] - tc;
                        p[269] = p[269] + tc;
                        p[273] = p[273] + tc;
                end
                256: begin
                        tc = f[255];
                        p[254] = p[254] - tc;
                        p[45] = p[45] + tc;
                end
                257: begin
                        tc = f[256];
                        p[45] = p[45] - tc;
                end
                258: begin
                        tc = f[257];
                        p[274] = p[274] - tc;
                        p[255] = p[255] + tc;
                end
                259: begin
                        tc = f[258];
                        p[8] = p[8] - tc;
                        p[274] = p[274] + tc;
                end
                260: begin
                        tc = f[259];
                        p[281] = p[281] - tc;
                        p[277] = p[277] + tc;
                end
                261: begin
                        tc = f[260];
                        p[275] = p[275] - tc;
                end
                262: begin
                        tc = f[261];
                        p[279] = p[279] - tc;
                        p[281] = p[281] + tc;
                end
                263: begin
                        tc = f[262];
                        p[276] = p[276] - tc*2;
                        p[282] = p[282] + tc;
                end
                264: begin
                        tc = f[263];
                        p[283] = p[283] - tc;
                        p[280] = p[280] + tc;
                end
                265: begin
                        tc = f[264];
                        p[276] = p[276] - tc;
                        p[285] = p[285] - tc;
                        p[284] = p[284] + tc;
                end
                266: begin
                        tc = f[265];
                        p[286] = p[286] - tc;
                        p[283] = p[283] + tc;
                end
                267: begin
                        tc = f[266];
                        p[275] = p[275] - tc;
                        p[278] = p[278] + tc;
                        p[287] = p[287] + tc;
                end
                268: begin
                        tc = f[267];
                        p[275] = p[275] - tc;
                        p[287] = p[287] + tc;
                end
                269: begin
                        tc = f[268];
                        p[288] = p[288] - tc;
                        p[286] = p[286] + tc;
                end
                270: begin
                        tc = f[269];
                        p[282] = p[282] - tc;
                        p[276] = p[276] + tc;
                end
                271: begin
                        tc = f[270];
                        p[289] = p[289] - tc;
                        p[288] = p[288] + tc;
                end
                272: begin
                        tc = f[271];
                        p[287] = p[287] - tc;
                        p[275] = p[275] + tc*2;
                end
                273: begin
                        tc = f[272];
                        p[277] = p[277] - tc;
                        p[284] = p[284] - tc;
                        p[285] = p[285] + tc;
                        p[289] = p[289] + tc;
                end
                274: begin
                        tc = f[273];
                        p[277] = p[277] - tc;
                        p[289] = p[289] + tc;
                end
                275: begin
                        tc = f[274];
                        p[45] = p[45] - tc;
                        p[275] = p[275] + tc;
                        p[290] = p[290] + tc;
                end
                276: begin
                        tc = f[275];
                        p[290] = p[290] - tc;
                        p[45] = p[45] + tc;
                end
                277: begin
                        tc = f[276];
                        p[292] = p[292] - tc;
                        p[291] = p[291] + tc;
                end
                278: begin
                        tc = f[277];
                        p[293] = p[293] - tc;
                        p[292] = p[292] + tc;
                end
                279: begin
                        tc = f[278];
                        p[46] = p[46] - tc;
                        p[276] = p[276] + tc;
                        p[294] = p[294] + tc;
                end
                280: begin
                        tc = f[279];
                        p[294] = p[294] - tc;
                        p[46] = p[46] + tc;
                end
                281: begin
                        tc = f[280];
                        p[296] = p[296] - tc;
                        p[295] = p[295] + tc;
                end
                282: begin
                        tc = f[281];
                        p[297] = p[297] - tc;
                        p[296] = p[296] + tc;
                end
                283: begin
                        tc = f[282];
                        p[291] = p[291] - tc;
                        p[295] = p[295] - tc;
                        p[8] = p[8] + tc;
                end
                284: begin
                        tc = f[283];
                        p[277] = p[277] - tc;
                        p[293] = p[293] + tc;
                        p[297] = p[297] + tc;
                end
                285: begin
                        tc = f[284];
                        p[278] = p[278] - tc;
                        p[47] = p[47] + tc;
                end
                286: begin
                        tc = f[285];
                        p[47] = p[47] - tc;
                end
                287: begin
                        tc = f[286];
                        p[298] = p[298] - tc;
                        p[279] = p[279] + tc;
                end
                288: begin
                        tc = f[287];
                        p[9] = p[9] - tc;
                        p[298] = p[298] + tc;
                end
                289: begin
                        tc = f[288];
                        p[305] = p[305] - tc;
                        p[301] = p[301] + tc;
                end
                290: begin
                        tc = f[289];
                        p[299] = p[299] - tc;
                end
                291: begin
                        tc = f[290];
                        p[303] = p[303] - tc;
                        p[305] = p[305] + tc;
                end
                292: begin
                        tc = f[291];
                        p[300] = p[300] - tc*2;
                        p[306] = p[306] + tc;
                end
                293: begin
                        tc = f[292];
                        p[307] = p[307] - tc;
                        p[304] = p[304] + tc;
                end
                294: begin
                        tc = f[293];
                        p[300] = p[300] - tc;
                        p[309] = p[309] - tc;
                        p[308] = p[308] + tc;
                end
                295: begin
                        tc = f[294];
                        p[310] = p[310] - tc;
                        p[307] = p[307] + tc;
                end
                296: begin
                        tc = f[295];
                        p[299] = p[299] - tc;
                        p[302] = p[302] + tc;
                        p[311] = p[311] + tc;
                end
                297: begin
                        tc = f[296];
                        p[299] = p[299] - tc;
                        p[311] = p[311] + tc;
                end
                298: begin
                        tc = f[297];
                        p[312] = p[312] - tc;
                        p[310] = p[310] + tc;
                end
                299: begin
                        tc = f[298];
                        p[306] = p[306] - tc;
                        p[300] = p[300] + tc;
                end
                300: begin
                        tc = f[299];
                        p[313] = p[313] - tc;
                        p[312] = p[312] + tc;
                end
                301: begin
                        tc = f[300];
                        p[311] = p[311] - tc;
                        p[299] = p[299] + tc*2;
                end
                302: begin
                        tc = f[301];
                        p[301] = p[301] - tc;
                        p[308] = p[308] - tc;
                        p[309] = p[309] + tc;
                        p[313] = p[313] + tc;
                end
                303: begin
                        tc = f[302];
                        p[301] = p[301] - tc;
                        p[313] = p[313] + tc;
                end
                304: begin
                        tc = f[303];
                        p[47] = p[47] - tc;
                        p[299] = p[299] + tc;
                        p[314] = p[314] + tc;
                end
                305: begin
                        tc = f[304];
                        p[314] = p[314] - tc;
                        p[47] = p[47] + tc;
                end
                306: begin
                        tc = f[305];
                        p[316] = p[316] - tc;
                        p[315] = p[315] + tc;
                end
                307: begin
                        tc = f[306];
                        p[317] = p[317] - tc;
                        p[316] = p[316] + tc;
                end
                308: begin
                        tc = f[307];
                        p[48] = p[48] - tc;
                        p[300] = p[300] + tc;
                        p[318] = p[318] + tc;
                end
                309: begin
                        tc = f[308];
                        p[318] = p[318] - tc;
                        p[48] = p[48] + tc;
                end
                310: begin
                        tc = f[309];
                        p[320] = p[320] - tc;
                        p[319] = p[319] + tc;
                end
                311: begin
                        tc = f[310];
                        p[321] = p[321] - tc;
                        p[320] = p[320] + tc;
                end
                312: begin
                        tc = f[311];
                        p[315] = p[315] - tc;
                        p[319] = p[319] - tc;
                        p[9] = p[9] + tc;
                end
                313: begin
                        tc = f[312];
                        p[301] = p[301] - tc;
                        p[317] = p[317] + tc;
                        p[321] = p[321] + tc;
                end
                314: begin
                        tc = f[313];
                        p[302] = p[302] - tc;
                        p[49] = p[49] + tc;
                end
                315: begin
                        tc = f[314];
                        p[49] = p[49] - tc;
                end
                316: begin
                        tc = f[315];
                        p[322] = p[322] - tc;
                        p[303] = p[303] + tc;
                end
                317: begin
                        tc = f[316];
                        p[10] = p[10] - tc;
                        p[322] = p[322] + tc;
                end
                318: begin
                        tc = f[317];
                        p[329] = p[329] - tc;
                        p[325] = p[325] + tc;
                end
                319: begin
                        tc = f[318];
                        p[323] = p[323] - tc;
                end
                320: begin
                        tc = f[319];
                        p[327] = p[327] - tc;
                        p[329] = p[329] + tc;
                end
                321: begin
                        tc = f[320];
                        p[324] = p[324] - tc*2;
                        p[330] = p[330] + tc;
                end
                322: begin
                        tc = f[321];
                        p[331] = p[331] - tc;
                        p[328] = p[328] + tc;
                end
                323: begin
                        tc = f[322];
                        p[324] = p[324] - tc;
                        p[333] = p[333] - tc;
                        p[332] = p[332] + tc;
                end
                324: begin
                        tc = f[323];
                        p[334] = p[334] - tc;
                        p[331] = p[331] + tc;
                end
                325: begin
                        tc = f[324];
                        p[323] = p[323] - tc;
                        p[326] = p[326] + tc;
                        p[335] = p[335] + tc;
                end
                326: begin
                        tc = f[325];
                        p[323] = p[323] - tc;
                        p[335] = p[335] + tc;
                end
                327: begin
                        tc = f[326];
                        p[336] = p[336] - tc;
                        p[334] = p[334] + tc;
                end
                328: begin
                        tc = f[327];
                        p[330] = p[330] - tc;
                        p[324] = p[324] + tc;
                end
                329: begin
                        tc = f[328];
                        p[337] = p[337] - tc;
                        p[336] = p[336] + tc;
                end
                330: begin
                        tc = f[329];
                        p[335] = p[335] - tc;
                        p[323] = p[323] + tc*2;
                end
                331: begin
                        tc = f[330];
                        p[325] = p[325] - tc;
                        p[332] = p[332] - tc;
                        p[333] = p[333] + tc;
                        p[337] = p[337] + tc;
                end
                332: begin
                        tc = f[331];
                        p[325] = p[325] - tc;
                        p[337] = p[337] + tc;
                end
                333: begin
                        tc = f[332];
                        p[49] = p[49] - tc;
                        p[323] = p[323] + tc;
                        p[338] = p[338] + tc;
                end
                334: begin
                        tc = f[333];
                        p[338] = p[338] - tc;
                        p[49] = p[49] + tc;
                end
                335: begin
                        tc = f[334];
                        p[340] = p[340] - tc;
                        p[339] = p[339] + tc;
                end
                336: begin
                        tc = f[335];
                        p[341] = p[341] - tc;
                        p[340] = p[340] + tc;
                end
                337: begin
                        tc = f[336];
                        p[50] = p[50] - tc;
                        p[324] = p[324] + tc;
                        p[342] = p[342] + tc;
                end
                338: begin
                        tc = f[337];
                        p[342] = p[342] - tc;
                        p[50] = p[50] + tc;
                end
                339: begin
                        tc = f[338];
                        p[344] = p[344] - tc;
                        p[343] = p[343] + tc;
                end
                340: begin
                        tc = f[339];
                        p[345] = p[345] - tc;
                        p[344] = p[344] + tc;
                end
                341: begin
                        tc = f[340];
                        p[339] = p[339] - tc;
                        p[343] = p[343] - tc;
                        p[10] = p[10] + tc;
                end
                342: begin
                        tc = f[341];
                        p[325] = p[325] - tc;
                        p[341] = p[341] + tc;
                        p[345] = p[345] + tc;
                end
                343: begin
                        tc = f[342];
                        p[326] = p[326] - tc;
                        p[51] = p[51] + tc;
                end
                344: begin
                        tc = f[343];
                        p[51] = p[51] - tc;
                end
                345: begin
                        tc = f[344];
                        p[346] = p[346] - tc;
                        p[327] = p[327] + tc;
                end
                346: begin
                        tc = f[345];
                        p[11] = p[11] - tc;
                        p[346] = p[346] + tc;
                end
                347: begin
                        tc = f[346];
                        p[348] = p[348] - tc;
                        p[349] = p[349] + tc;
                end
                348: begin
                        tc = f[347];
                        p[351] = p[351] - tc;
                        p[350] = p[350] + tc;
                end
                349: begin
                        tc = f[348];
                        p[40] = p[40] - tc;
                        p[347] = p[347] + tc;
                        p[352] = p[352] + tc;
                end
                350: begin
                        tc = f[349];
                        p[352] = p[352] - tc;
                        p[40] = p[40] + tc;
                end
                351: begin
                        tc = f[350];
                        p[354] = p[354] - tc;
                        p[353] = p[353] + tc;
                end
                352: begin
                        tc = f[351];
                        p[355] = p[355] - tc;
                        p[354] = p[354] + tc;
                end
                353: begin
                        tc = f[352];
                        p[51] = p[51] - tc;
                        p[348] = p[348] + tc;
                        p[356] = p[356] + tc;
                end
                354: begin
                        tc = f[353];
                        p[356] = p[356] - tc;
                        p[51] = p[51] + tc;
                end
                355: begin
                        tc = f[354];
                        p[358] = p[358] - tc;
                        p[357] = p[357] + tc;
                end
                356: begin
                        tc = f[355];
                        p[359] = p[359] - tc;
                        p[358] = p[358] + tc;
                end
                357: begin
                        tc = f[356];
                        p[353] = p[353] - tc;
                        p[357] = p[357] - tc;
                        p[11] = p[11] + tc;
                end
                358: begin
                        tc = f[357];
                        p[350] = p[350] - tc;
                        p[355] = p[355] + tc;
                        p[359] = p[359] + tc;
                end
                359: begin
                        tc = f[358];
                        p[349] = p[349] - tc;
                        p[52] = p[52] + tc;
                end
                360: begin
                        tc = f[359];
                        p[52] = p[52] - tc;
                end
                361: begin
                        tc = f[360];
                        p[360] = p[360] - tc;
                        p[351] = p[351] + tc;
                end
                362: begin
                        tc = f[361];
                        p[12] = p[12] - tc;
                        p[360] = p[360] + tc;
                end
                363: begin
                        tc = f[362];
                        p[367] = p[367] - tc;
                        p[363] = p[363] + tc;
                end
                364: begin
                        tc = f[363];
                        p[361] = p[361] - tc;
                end
                365: begin
                        tc = f[364];
                        p[365] = p[365] - tc;
                        p[367] = p[367] + tc;
                end
                366: begin
                        tc = f[365];
                        p[362] = p[362] - tc*2;
                        p[368] = p[368] + tc;
                end
                367: begin
                        tc = f[366];
                        p[369] = p[369] - tc;
                        p[366] = p[366] + tc;
                end
                368: begin
                        tc = f[367];
                        p[362] = p[362] - tc;
                        p[371] = p[371] - tc;
                        p[370] = p[370] + tc;
                end
                369: begin
                        tc = f[368];
                        p[372] = p[372] - tc;
                        p[369] = p[369] + tc;
                end
                370: begin
                        tc = f[369];
                        p[361] = p[361] - tc;
                        p[364] = p[364] + tc;
                        p[373] = p[373] + tc;
                end
                371: begin
                        tc = f[370];
                        p[361] = p[361] - tc;
                        p[373] = p[373] + tc;
                end
                372: begin
                        tc = f[371];
                        p[374] = p[374] - tc;
                        p[372] = p[372] + tc;
                end
                373: begin
                        tc = f[372];
                        p[368] = p[368] - tc;
                        p[362] = p[362] + tc;
                end
                374: begin
                        tc = f[373];
                        p[375] = p[375] - tc;
                        p[374] = p[374] + tc;
                end
                375: begin
                        tc = f[374];
                        p[373] = p[373] - tc;
                        p[361] = p[361] + tc*2;
                end
                376: begin
                        tc = f[375];
                        p[363] = p[363] - tc;
                        p[370] = p[370] - tc;
                        p[371] = p[371] + tc;
                        p[375] = p[375] + tc;
                end
                377: begin
                        tc = f[376];
                        p[363] = p[363] - tc;
                        p[375] = p[375] + tc;
                end
                378: begin
                        tc = f[377];
                        p[53] = p[53] - tc;
                        p[361] = p[361] + tc;
                        p[376] = p[376] + tc;
                end
                379: begin
                        tc = f[378];
                        p[376] = p[376] - tc;
                        p[53] = p[53] + tc;
                end
                380: begin
                        tc = f[379];
                        p[378] = p[378] - tc;
                        p[377] = p[377] + tc;
                end
                381: begin
                        tc = f[380];
                        p[379] = p[379] - tc;
                        p[378] = p[378] + tc;
                end
                382: begin
                        tc = f[381];
                        p[54] = p[54] - tc;
                        p[362] = p[362] + tc;
                        p[380] = p[380] + tc;
                end
                383: begin
                        tc = f[382];
                        p[380] = p[380] - tc;
                        p[54] = p[54] + tc;
                end
                384: begin
                        tc = f[383];
                        p[382] = p[382] - tc;
                        p[381] = p[381] + tc;
                end
                385: begin
                        tc = f[384];
                        p[383] = p[383] - tc;
                        p[382] = p[382] + tc;
                end
                386: begin
                        tc = f[385];
                        p[377] = p[377] - tc;
                        p[381] = p[381] - tc;
                        p[12] = p[12] + tc;
                end
                387: begin
                        tc = f[386];
                        p[363] = p[363] - tc;
                        p[379] = p[379] + tc;
                        p[383] = p[383] + tc;
                end
                388: begin
                        tc = f[387];
                        p[364] = p[364] - tc;
                        p[55] = p[55] + tc;
                end
                389: begin
                        tc = f[388];
                        p[55] = p[55] - tc;
                end
                390: begin
                        tc = f[389];
                        p[384] = p[384] - tc;
                        p[365] = p[365] + tc;
                end
                391: begin
                        tc = f[390];
                        p[13] = p[13] - tc;
                        p[384] = p[384] + tc;
                end
                392: begin
                        tc = f[391];
                        p[391] = p[391] - tc;
                        p[387] = p[387] + tc;
                end
                393: begin
                        tc = f[392];
                        p[385] = p[385] - tc;
                end
                394: begin
                        tc = f[393];
                        p[389] = p[389] - tc;
                        p[391] = p[391] + tc;
                end
                395: begin
                        tc = f[394];
                        p[386] = p[386] - tc*2;
                        p[392] = p[392] + tc;
                end
                396: begin
                        tc = f[395];
                        p[393] = p[393] - tc;
                        p[390] = p[390] + tc;
                end
                397: begin
                        tc = f[396];
                        p[386] = p[386] - tc;
                        p[395] = p[395] - tc;
                        p[394] = p[394] + tc;
                end
                398: begin
                        tc = f[397];
                        p[396] = p[396] - tc;
                        p[393] = p[393] + tc;
                end
                399: begin
                        tc = f[398];
                        p[385] = p[385] - tc;
                        p[388] = p[388] + tc;
                        p[397] = p[397] + tc;
                end
                400: begin
                        tc = f[399];
                        p[385] = p[385] - tc;
                        p[397] = p[397] + tc;
                end
                401: begin
                        tc = f[400];
                        p[398] = p[398] - tc;
                        p[396] = p[396] + tc;
                end
                402: begin
                        tc = f[401];
                        p[392] = p[392] - tc;
                        p[386] = p[386] + tc;
                end
                403: begin
                        tc = f[402];
                        p[399] = p[399] - tc;
                        p[398] = p[398] + tc;
                end
                404: begin
                        tc = f[403];
                        p[397] = p[397] - tc;
                        p[385] = p[385] + tc*2;
                end
                405: begin
                        tc = f[404];
                        p[387] = p[387] - tc;
                        p[394] = p[394] - tc;
                        p[395] = p[395] + tc;
                        p[399] = p[399] + tc;
                end
                406: begin
                        tc = f[405];
                        p[387] = p[387] - tc;
                        p[399] = p[399] + tc;
                end
                407: begin
                        tc = f[406];
                        p[55] = p[55] - tc;
                        p[385] = p[385] + tc;
                        p[400] = p[400] + tc;
                end
                408: begin
                        tc = f[407];
                        p[400] = p[400] - tc;
                        p[55] = p[55] + tc;
                end
                409: begin
                        tc = f[408];
                        p[402] = p[402] - tc;
                        p[401] = p[401] + tc;
                end
                410: begin
                        tc = f[409];
                        p[403] = p[403] - tc;
                        p[402] = p[402] + tc;
                end
                411: begin
                        tc = f[410];
                        p[56] = p[56] - tc;
                        p[386] = p[386] + tc;
                        p[404] = p[404] + tc;
                end
                412: begin
                        tc = f[411];
                        p[404] = p[404] - tc;
                        p[56] = p[56] + tc;
                end
                413: begin
                        tc = f[412];
                        p[406] = p[406] - tc;
                        p[405] = p[405] + tc;
                end
                414: begin
                        tc = f[413];
                        p[407] = p[407] - tc;
                        p[406] = p[406] + tc;
                end
                415: begin
                        tc = f[414];
                        p[401] = p[401] - tc;
                        p[405] = p[405] - tc;
                        p[13] = p[13] + tc;
                end
                416: begin
                        tc = f[415];
                        p[387] = p[387] - tc;
                        p[403] = p[403] + tc;
                        p[407] = p[407] + tc;
                end
                417: begin
                        tc = f[416];
                        p[388] = p[388] - tc;
                        p[57] = p[57] + tc;
                end
                418: begin
                        tc = f[417];
                        p[57] = p[57] - tc;
                end
                419: begin
                        tc = f[418];
                        p[408] = p[408] - tc;
                        p[389] = p[389] + tc;
                end
                420: begin
                        tc = f[419];
                        p[14] = p[14] - tc;
                        p[408] = p[408] + tc;
                end
                421: begin
                        tc = f[420];
                        p[415] = p[415] - tc;
                        p[411] = p[411] + tc;
                end
                422: begin
                        tc = f[421];
                        p[409] = p[409] - tc;
                end
                423: begin
                        tc = f[422];
                        p[413] = p[413] - tc;
                        p[415] = p[415] + tc;
                end
                424: begin
                        tc = f[423];
                        p[410] = p[410] - tc*2;
                        p[416] = p[416] + tc;
                end
                425: begin
                        tc = f[424];
                        p[417] = p[417] - tc;
                        p[414] = p[414] + tc;
                end
                426: begin
                        tc = f[425];
                        p[410] = p[410] - tc;
                        p[419] = p[419] - tc;
                        p[418] = p[418] + tc;
                end
                427: begin
                        tc = f[426];
                        p[420] = p[420] - tc;
                        p[417] = p[417] + tc;
                end
                428: begin
                        tc = f[427];
                        p[409] = p[409] - tc;
                        p[412] = p[412] + tc;
                        p[421] = p[421] + tc;
                end
                429: begin
                        tc = f[428];
                        p[409] = p[409] - tc;
                        p[421] = p[421] + tc;
                end
                430: begin
                        tc = f[429];
                        p[422] = p[422] - tc;
                        p[420] = p[420] + tc;
                end
                431: begin
                        tc = f[430];
                        p[416] = p[416] - tc;
                        p[410] = p[410] + tc;
                end
                432: begin
                        tc = f[431];
                        p[423] = p[423] - tc;
                        p[422] = p[422] + tc;
                end
                433: begin
                        tc = f[432];
                        p[421] = p[421] - tc;
                        p[409] = p[409] + tc*2;
                end
                434: begin
                        tc = f[433];
                        p[411] = p[411] - tc;
                        p[418] = p[418] - tc;
                        p[419] = p[419] + tc;
                        p[423] = p[423] + tc;
                end
                435: begin
                        tc = f[434];
                        p[411] = p[411] - tc;
                        p[423] = p[423] + tc;
                end
                436: begin
                        tc = f[435];
                        p[57] = p[57] - tc;
                        p[409] = p[409] + tc;
                        p[424] = p[424] + tc;
                end
                437: begin
                        tc = f[436];
                        p[424] = p[424] - tc;
                        p[57] = p[57] + tc;
                end
                438: begin
                        tc = f[437];
                        p[426] = p[426] - tc;
                        p[425] = p[425] + tc;
                end
                439: begin
                        tc = f[438];
                        p[427] = p[427] - tc;
                        p[426] = p[426] + tc;
                end
                440: begin
                        tc = f[439];
                        p[58] = p[58] - tc;
                        p[410] = p[410] + tc;
                        p[428] = p[428] + tc;
                end
                441: begin
                        tc = f[440];
                        p[428] = p[428] - tc;
                        p[58] = p[58] + tc;
                end
                442: begin
                        tc = f[441];
                        p[430] = p[430] - tc;
                        p[429] = p[429] + tc;
                end
                443: begin
                        tc = f[442];
                        p[431] = p[431] - tc;
                        p[430] = p[430] + tc;
                end
                444: begin
                        tc = f[443];
                        p[425] = p[425] - tc;
                        p[429] = p[429] - tc;
                        p[14] = p[14] + tc;
                end
                445: begin
                        tc = f[444];
                        p[411] = p[411] - tc;
                        p[427] = p[427] + tc;
                        p[431] = p[431] + tc;
                end
                446: begin
                        tc = f[445];
                        p[412] = p[412] - tc;
                        p[59] = p[59] + tc;
                end
                447: begin
                        tc = f[446];
                        p[59] = p[59] - tc;
                end
                448: begin
                        tc = f[447];
                        p[432] = p[432] - tc;
                        p[413] = p[413] + tc;
                end
                449: begin
                        tc = f[448];
                        p[15] = p[15] - tc;
                        p[432] = p[432] + tc;
                end
                450: begin
                        tc = f[449];
                        p[439] = p[439] - tc;
                        p[435] = p[435] + tc;
                end
                451: begin
                        tc = f[450];
                        p[433] = p[433] - tc;
                end
                452: begin
                        tc = f[451];
                        p[437] = p[437] - tc;
                        p[439] = p[439] + tc;
                end
                453: begin
                        tc = f[452];
                        p[434] = p[434] - tc*2;
                        p[440] = p[440] + tc;
                end
                454: begin
                        tc = f[453];
                        p[441] = p[441] - tc;
                        p[438] = p[438] + tc;
                end
                455: begin
                        tc = f[454];
                        p[434] = p[434] - tc;
                        p[443] = p[443] - tc;
                        p[442] = p[442] + tc;
                end
                456: begin
                        tc = f[455];
                        p[444] = p[444] - tc;
                        p[441] = p[441] + tc;
                end
                457: begin
                        tc = f[456];
                        p[433] = p[433] - tc;
                        p[436] = p[436] + tc;
                        p[445] = p[445] + tc;
                end
                458: begin
                        tc = f[457];
                        p[433] = p[433] - tc;
                        p[445] = p[445] + tc;
                end
                459: begin
                        tc = f[458];
                        p[446] = p[446] - tc;
                        p[444] = p[444] + tc;
                end
                460: begin
                        tc = f[459];
                        p[440] = p[440] - tc;
                        p[434] = p[434] + tc;
                end
                461: begin
                        tc = f[460];
                        p[447] = p[447] - tc;
                        p[446] = p[446] + tc;
                end
                462: begin
                        tc = f[461];
                        p[445] = p[445] - tc;
                        p[433] = p[433] + tc*2;
                end
                463: begin
                        tc = f[462];
                        p[435] = p[435] - tc;
                        p[442] = p[442] - tc;
                        p[443] = p[443] + tc;
                        p[447] = p[447] + tc;
                end
                464: begin
                        tc = f[463];
                        p[435] = p[435] - tc;
                        p[447] = p[447] + tc;
                end
                465: begin
                        tc = f[464];
                        p[59] = p[59] - tc;
                        p[433] = p[433] + tc;
                        p[448] = p[448] + tc;
                end
                466: begin
                        tc = f[465];
                        p[448] = p[448] - tc;
                        p[59] = p[59] + tc;
                end
                467: begin
                        tc = f[466];
                        p[450] = p[450] - tc;
                        p[449] = p[449] + tc;
                end
                468: begin
                        tc = f[467];
                        p[451] = p[451] - tc;
                        p[450] = p[450] + tc;
                end
                469: begin
                        tc = f[468];
                        p[60] = p[60] - tc;
                        p[434] = p[434] + tc;
                        p[452] = p[452] + tc;
                end
                470: begin
                        tc = f[469];
                        p[452] = p[452] - tc;
                        p[60] = p[60] + tc;
                end
                471: begin
                        tc = f[470];
                        p[454] = p[454] - tc;
                        p[453] = p[453] + tc;
                end
                472: begin
                        tc = f[471];
                        p[455] = p[455] - tc;
                        p[454] = p[454] + tc;
                end
                473: begin
                        tc = f[472];
                        p[449] = p[449] - tc;
                        p[453] = p[453] - tc;
                        p[15] = p[15] + tc;
                end
                474: begin
                        tc = f[473];
                        p[435] = p[435] - tc;
                        p[451] = p[451] + tc;
                        p[455] = p[455] + tc;
                end
                475: begin
                        tc = f[474];
                        p[436] = p[436] - tc;
                        p[61] = p[61] + tc;
                end
                476: begin
                        tc = f[475];
                        p[61] = p[61] - tc;
                end
                477: begin
                        tc = f[476];
                        p[456] = p[456] - tc;
                        p[437] = p[437] + tc;
                end
                478: begin
                        tc = f[477];
                        p[16] = p[16] - tc;
                        p[456] = p[456] + tc;
                end
                479: begin
                        tc = f[478];
                        p[458] = p[458] - tc;
                        p[459] = p[459] + tc;
                end
                480: begin
                        tc = f[479];
                        p[461] = p[461] - tc;
                        p[460] = p[460] + tc;
                end
                481: begin
                        tc = f[480];
                        p[61] = p[61] - tc;
                        p[457] = p[457] + tc;
                        p[462] = p[462] + tc;
                end
                482: begin
                        tc = f[481];
                        p[462] = p[462] - tc;
                        p[61] = p[61] + tc;
                end
                483: begin
                        tc = f[482];
                        p[464] = p[464] - tc;
                        p[463] = p[463] + tc;
                end
                484: begin
                        tc = f[483];
                        p[465] = p[465] - tc;
                        p[464] = p[464] + tc;
                end
                485: begin
                        tc = f[484];
                        p[52] = p[52] - tc;
                        p[458] = p[458] + tc;
                        p[466] = p[466] + tc;
                end
                486: begin
                        tc = f[485];
                        p[466] = p[466] - tc;
                        p[52] = p[52] + tc;
                end
                487: begin
                        tc = f[486];
                        p[468] = p[468] - tc;
                        p[467] = p[467] + tc;
                end
                488: begin
                        tc = f[487];
                        p[469] = p[469] - tc;
                        p[468] = p[468] + tc;
                end
                489: begin
                        tc = f[488];
                        p[463] = p[463] - tc;
                        p[467] = p[467] - tc;
                        p[16] = p[16] + tc;
                end
                490: begin
                        tc = f[489];
                        p[460] = p[460] - tc;
                        p[465] = p[465] + tc;
                        p[469] = p[469] + tc;
                end
                491: begin
                        tc = f[490];
                        p[459] = p[459] - tc;
                        p[62] = p[62] + tc;
                end
                492: begin
                        tc = f[491];
                        p[62] = p[62] - tc;
                end
                493: begin
                        tc = f[492];
                        p[470] = p[470] - tc;
                        p[461] = p[461] + tc;
                end
                494: begin
                        tc = f[493];
                        p[17] = p[17] - tc;
                        p[470] = p[470] + tc;
                end
                495: begin
                        tc = f[494];
                        p[477] = p[477] - tc;
                        p[473] = p[473] + tc;
                end
                496: begin
                        tc = f[495];
                        p[471] = p[471] - tc;
                end
                497: begin
                        tc = f[496];
                        p[475] = p[475] - tc;
                        p[477] = p[477] + tc;
                end
                498: begin
                        tc = f[497];
                        p[472] = p[472] - tc*2;
                        p[478] = p[478] + tc;
                end
                499: begin
                        tc = f[498];
                        p[479] = p[479] - tc;
                        p[476] = p[476] + tc;
                end
                500: begin
                        tc = f[499];
                        p[472] = p[472] - tc;
                        p[481] = p[481] - tc;
                        p[480] = p[480] + tc;
                end
                501: begin
                        tc = f[500];
                        p[482] = p[482] - tc;
                        p[479] = p[479] + tc;
                end
                502: begin
                        tc = f[501];
                        p[471] = p[471] - tc;
                        p[474] = p[474] + tc;
                        p[483] = p[483] + tc;
                end
                503: begin
                        tc = f[502];
                        p[471] = p[471] - tc;
                        p[483] = p[483] + tc;
                end
                504: begin
                        tc = f[503];
                        p[484] = p[484] - tc;
                        p[482] = p[482] + tc;
                end
                505: begin
                        tc = f[504];
                        p[478] = p[478] - tc;
                        p[472] = p[472] + tc;
                end
                506: begin
                        tc = f[505];
                        p[485] = p[485] - tc;
                        p[484] = p[484] + tc;
                end
                507: begin
                        tc = f[506];
                        p[483] = p[483] - tc;
                        p[471] = p[471] + tc*2;
                end
                508: begin
                        tc = f[507];
                        p[473] = p[473] - tc;
                        p[480] = p[480] - tc;
                        p[481] = p[481] + tc;
                        p[485] = p[485] + tc;
                end
                509: begin
                        tc = f[508];
                        p[473] = p[473] - tc;
                        p[485] = p[485] + tc;
                end
                510: begin
                        tc = f[509];
                        p[63] = p[63] - tc;
                        p[471] = p[471] + tc;
                        p[486] = p[486] + tc;
                end
                511: begin
                        tc = f[510];
                        p[486] = p[486] - tc;
                        p[63] = p[63] + tc;
                end
                512: begin
                        tc = f[511];
                        p[488] = p[488] - tc;
                        p[487] = p[487] + tc;
                end
                513: begin
                        tc = f[512];
                        p[489] = p[489] - tc;
                        p[488] = p[488] + tc;
                end
                514: begin
                        tc = f[513];
                        p[64] = p[64] - tc;
                        p[472] = p[472] + tc;
                        p[490] = p[490] + tc;
                end
                515: begin
                        tc = f[514];
                        p[490] = p[490] - tc;
                        p[64] = p[64] + tc;
                end
                516: begin
                        tc = f[515];
                        p[492] = p[492] - tc;
                        p[491] = p[491] + tc;
                end
                517: begin
                        tc = f[516];
                        p[493] = p[493] - tc;
                        p[492] = p[492] + tc;
                end
                518: begin
                        tc = f[517];
                        p[487] = p[487] - tc;
                        p[491] = p[491] - tc;
                        p[17] = p[17] + tc;
                end
                519: begin
                        tc = f[518];
                        p[473] = p[473] - tc;
                        p[489] = p[489] + tc;
                        p[493] = p[493] + tc;
                end
                520: begin
                        tc = f[519];
                        p[474] = p[474] - tc;
                        p[65] = p[65] + tc;
                end
                521: begin
                        tc = f[520];
                        p[65] = p[65] - tc;
                end
                522: begin
                        tc = f[521];
                        p[494] = p[494] - tc;
                        p[475] = p[475] + tc;
                end
                523: begin
                        tc = f[522];
                        p[18] = p[18] - tc;
                        p[494] = p[494] + tc;
                end
                524: begin
                        tc = f[523];
                        p[501] = p[501] - tc;
                        p[497] = p[497] + tc;
                end
                525: begin
                        tc = f[524];
                        p[495] = p[495] - tc;
                end
                526: begin
                        tc = f[525];
                        p[499] = p[499] - tc;
                        p[501] = p[501] + tc;
                end
                527: begin
                        tc = f[526];
                        p[496] = p[496] - tc*2;
                        p[502] = p[502] + tc;
                end
                528: begin
                        tc = f[527];
                        p[503] = p[503] - tc;
                        p[500] = p[500] + tc;
                end
                529: begin
                        tc = f[528];
                        p[496] = p[496] - tc;
                        p[505] = p[505] - tc;
                        p[504] = p[504] + tc;
                end
                530: begin
                        tc = f[529];
                        p[506] = p[506] - tc;
                        p[503] = p[503] + tc;
                end
                531: begin
                        tc = f[530];
                        p[495] = p[495] - tc;
                        p[498] = p[498] + tc;
                        p[507] = p[507] + tc;
                end
                532: begin
                        tc = f[531];
                        p[495] = p[495] - tc;
                        p[507] = p[507] + tc;
                end
                533: begin
                        tc = f[532];
                        p[508] = p[508] - tc;
                        p[506] = p[506] + tc;
                end
                534: begin
                        tc = f[533];
                        p[502] = p[502] - tc;
                        p[496] = p[496] + tc;
                end
                535: begin
                        tc = f[534];
                        p[509] = p[509] - tc;
                        p[508] = p[508] + tc;
                end
                536: begin
                        tc = f[535];
                        p[507] = p[507] - tc;
                        p[495] = p[495] + tc*2;
                end
                537: begin
                        tc = f[536];
                        p[497] = p[497] - tc;
                        p[504] = p[504] - tc;
                        p[505] = p[505] + tc;
                        p[509] = p[509] + tc;
                end
                538: begin
                        tc = f[537];
                        p[497] = p[497] - tc;
                        p[509] = p[509] + tc;
                end
                539: begin
                        tc = f[538];
                        p[65] = p[65] - tc;
                        p[495] = p[495] + tc;
                        p[510] = p[510] + tc;
                end
                540: begin
                        tc = f[539];
                        p[510] = p[510] - tc;
                        p[65] = p[65] + tc;
                end
                541: begin
                        tc = f[540];
                        p[512] = p[512] - tc;
                        p[511] = p[511] + tc;
                end
                542: begin
                        tc = f[541];
                        p[513] = p[513] - tc;
                        p[512] = p[512] + tc;
                end
                543: begin
                        tc = f[542];
                        p[66] = p[66] - tc;
                        p[496] = p[496] + tc;
                        p[514] = p[514] + tc;
                end
                544: begin
                        tc = f[543];
                        p[514] = p[514] - tc;
                        p[66] = p[66] + tc;
                end
                545: begin
                        tc = f[544];
                        p[516] = p[516] - tc;
                        p[515] = p[515] + tc;
                end
                546: begin
                        tc = f[545];
                        p[517] = p[517] - tc;
                        p[516] = p[516] + tc;
                end
                547: begin
                        tc = f[546];
                        p[511] = p[511] - tc;
                        p[515] = p[515] - tc;
                        p[18] = p[18] + tc;
                end
                548: begin
                        tc = f[547];
                        p[497] = p[497] - tc;
                        p[513] = p[513] + tc;
                        p[517] = p[517] + tc;
                end
                549: begin
                        tc = f[548];
                        p[498] = p[498] - tc;
                        p[67] = p[67] + tc;
                end
                550: begin
                        tc = f[549];
                        p[67] = p[67] - tc;
                end
                551: begin
                        tc = f[550];
                        p[518] = p[518] - tc;
                        p[499] = p[499] + tc;
                end
                552: begin
                        tc = f[551];
                        p[19] = p[19] - tc;
                        p[518] = p[518] + tc;
                end
                553: begin
                        tc = f[552];
                        p[525] = p[525] - tc;
                        p[521] = p[521] + tc;
                end
                554: begin
                        tc = f[553];
                        p[519] = p[519] - tc;
                end
                555: begin
                        tc = f[554];
                        p[523] = p[523] - tc;
                        p[525] = p[525] + tc;
                end
                556: begin
                        tc = f[555];
                        p[520] = p[520] - tc*2;
                        p[526] = p[526] + tc;
                end
                557: begin
                        tc = f[556];
                        p[527] = p[527] - tc;
                        p[524] = p[524] + tc;
                end
                558: begin
                        tc = f[557];
                        p[520] = p[520] - tc;
                        p[529] = p[529] - tc;
                        p[528] = p[528] + tc;
                end
                559: begin
                        tc = f[558];
                        p[530] = p[530] - tc;
                        p[527] = p[527] + tc;
                end
                560: begin
                        tc = f[559];
                        p[519] = p[519] - tc;
                        p[522] = p[522] + tc;
                        p[531] = p[531] + tc;
                end
                561: begin
                        tc = f[560];
                        p[519] = p[519] - tc;
                        p[531] = p[531] + tc;
                end
                562: begin
                        tc = f[561];
                        p[532] = p[532] - tc;
                        p[530] = p[530] + tc;
                end
                563: begin
                        tc = f[562];
                        p[526] = p[526] - tc;
                        p[520] = p[520] + tc;
                end
                564: begin
                        tc = f[563];
                        p[533] = p[533] - tc;
                        p[532] = p[532] + tc;
                end
                565: begin
                        tc = f[564];
                        p[531] = p[531] - tc;
                        p[519] = p[519] + tc*2;
                end
                566: begin
                        tc = f[565];
                        p[521] = p[521] - tc;
                        p[528] = p[528] - tc;
                        p[529] = p[529] + tc;
                        p[533] = p[533] + tc;
                end
                567: begin
                        tc = f[566];
                        p[521] = p[521] - tc;
                        p[533] = p[533] + tc;
                end
                568: begin
                        tc = f[567];
                        p[67] = p[67] - tc;
                        p[519] = p[519] + tc;
                        p[534] = p[534] + tc;
                end
                569: begin
                        tc = f[568];
                        p[534] = p[534] - tc;
                        p[67] = p[67] + tc;
                end
                570: begin
                        tc = f[569];
                        p[536] = p[536] - tc;
                        p[535] = p[535] + tc;
                end
                571: begin
                        tc = f[570];
                        p[537] = p[537] - tc;
                        p[536] = p[536] + tc;
                end
                572: begin
                        tc = f[571];
                        p[68] = p[68] - tc;
                        p[520] = p[520] + tc;
                        p[538] = p[538] + tc;
                end
                573: begin
                        tc = f[572];
                        p[538] = p[538] - tc;
                        p[68] = p[68] + tc;
                end
                574: begin
                        tc = f[573];
                        p[540] = p[540] - tc;
                        p[539] = p[539] + tc;
                end
                575: begin
                        tc = f[574];
                        p[541] = p[541] - tc;
                        p[540] = p[540] + tc;
                end
                576: begin
                        tc = f[575];
                        p[535] = p[535] - tc;
                        p[539] = p[539] - tc;
                        p[19] = p[19] + tc;
                end
                577: begin
                        tc = f[576];
                        p[521] = p[521] - tc;
                        p[537] = p[537] + tc;
                        p[541] = p[541] + tc;
                end
                578: begin
                        tc = f[577];
                        p[522] = p[522] - tc;
                        p[69] = p[69] + tc;
                end
                579: begin
                        tc = f[578];
                        p[69] = p[69] - tc;
                end
                580: begin
                        tc = f[579];
                        p[542] = p[542] - tc;
                        p[523] = p[523] + tc;
                end
                581: begin
                        tc = f[580];
                        p[20] = p[20] - tc;
                        p[542] = p[542] + tc;
                end
                582: begin
                        tc = f[581];
                        p[544] = p[544] - tc;
                        p[545] = p[545] + tc;
                end
                583: begin
                        tc = f[582];
                        p[547] = p[547] - tc;
                        p[546] = p[546] + tc;
                end
                584: begin
                        tc = f[583];
                        p[69] = p[69] - tc;
                        p[543] = p[543] + tc;
                        p[548] = p[548] + tc;
                end
                585: begin
                        tc = f[584];
                        p[548] = p[548] - tc;
                        p[69] = p[69] + tc;
                end
                586: begin
                        tc = f[585];
                        p[550] = p[550] - tc;
                        p[549] = p[549] + tc;
                end
                587: begin
                        tc = f[586];
                        p[551] = p[551] - tc;
                        p[550] = p[550] + tc;
                end
                588: begin
                        tc = f[587];
                        p[62] = p[62] - tc;
                        p[544] = p[544] + tc;
                        p[552] = p[552] + tc;
                end
                589: begin
                        tc = f[588];
                        p[552] = p[552] - tc;
                        p[62] = p[62] + tc;
                end
                590: begin
                        tc = f[589];
                        p[554] = p[554] - tc;
                        p[553] = p[553] + tc;
                end
                591: begin
                        tc = f[590];
                        p[555] = p[555] - tc;
                        p[554] = p[554] + tc;
                end
                592: begin
                        tc = f[591];
                        p[549] = p[549] - tc;
                        p[553] = p[553] - tc;
                        p[20] = p[20] + tc;
                end
                593: begin
                        tc = f[592];
                        p[546] = p[546] - tc;
                        p[551] = p[551] + tc;
                        p[555] = p[555] + tc;
                end
                594: begin
                        tc = f[593];
                        p[545] = p[545] - tc;
                        p[70] = p[70] + tc;
                end
                595: begin
                        tc = f[594];
                        p[70] = p[70] - tc;
                end
                596: begin
                        tc = f[595];
                        p[556] = p[556] - tc;
                        p[547] = p[547] + tc;
                end
                597: begin
                        tc = f[596];
                        p[21] = p[21] - tc;
                        p[556] = p[556] + tc;
                end
                598: begin
                        tc = f[597];
                        p[563] = p[563] - tc;
                        p[559] = p[559] + tc;
                end
                599: begin
                        tc = f[598];
                        p[557] = p[557] - tc;
                end
                600: begin
                        tc = f[599];
                        p[561] = p[561] - tc;
                        p[563] = p[563] + tc;
                end
                601: begin
                        tc = f[600];
                        p[558] = p[558] - tc*2;
                        p[564] = p[564] + tc;
                end
                602: begin
                        tc = f[601];
                        p[565] = p[565] - tc;
                        p[562] = p[562] + tc;
                end
                603: begin
                        tc = f[602];
                        p[558] = p[558] - tc;
                        p[567] = p[567] - tc;
                        p[566] = p[566] + tc;
                end
                604: begin
                        tc = f[603];
                        p[568] = p[568] - tc;
                        p[565] = p[565] + tc;
                end
                605: begin
                        tc = f[604];
                        p[557] = p[557] - tc;
                        p[560] = p[560] + tc;
                        p[569] = p[569] + tc;
                end
                606: begin
                        tc = f[605];
                        p[557] = p[557] - tc;
                        p[569] = p[569] + tc;
                end
                607: begin
                        tc = f[606];
                        p[570] = p[570] - tc;
                        p[568] = p[568] + tc;
                end
                608: begin
                        tc = f[607];
                        p[564] = p[564] - tc;
                        p[558] = p[558] + tc;
                end
                609: begin
                        tc = f[608];
                        p[571] = p[571] - tc;
                        p[570] = p[570] + tc;
                end
                610: begin
                        tc = f[609];
                        p[569] = p[569] - tc;
                        p[557] = p[557] + tc*2;
                end
                611: begin
                        tc = f[610];
                        p[559] = p[559] - tc;
                        p[566] = p[566] - tc;
                        p[567] = p[567] + tc;
                        p[571] = p[571] + tc;
                end
                612: begin
                        tc = f[611];
                        p[559] = p[559] - tc;
                        p[571] = p[571] + tc;
                end
                613: begin
                        tc = f[612];
                        p[71] = p[71] - tc;
                        p[557] = p[557] + tc;
                        p[572] = p[572] + tc;
                end
                614: begin
                        tc = f[613];
                        p[572] = p[572] - tc;
                        p[71] = p[71] + tc;
                end
                615: begin
                        tc = f[614];
                        p[574] = p[574] - tc;
                        p[573] = p[573] + tc;
                end
                616: begin
                        tc = f[615];
                        p[575] = p[575] - tc;
                        p[574] = p[574] + tc;
                end
                617: begin
                        tc = f[616];
                        p[72] = p[72] - tc;
                        p[558] = p[558] + tc;
                        p[576] = p[576] + tc;
                end
                618: begin
                        tc = f[617];
                        p[576] = p[576] - tc;
                        p[72] = p[72] + tc;
                end
                619: begin
                        tc = f[618];
                        p[578] = p[578] - tc;
                        p[577] = p[577] + tc;
                end
                620: begin
                        tc = f[619];
                        p[579] = p[579] - tc;
                        p[578] = p[578] + tc;
                end
                621: begin
                        tc = f[620];
                        p[573] = p[573] - tc;
                        p[577] = p[577] - tc;
                        p[21] = p[21] + tc;
                end
                622: begin
                        tc = f[621];
                        p[559] = p[559] - tc;
                        p[575] = p[575] + tc;
                        p[579] = p[579] + tc;
                end
                623: begin
                        tc = f[622];
                        p[560] = p[560] - tc;
                        p[73] = p[73] + tc;
                end
                624: begin
                        tc = f[623];
                        p[73] = p[73] - tc;
                end
                625: begin
                        tc = f[624];
                        p[580] = p[580] - tc;
                        p[561] = p[561] + tc;
                end
                626: begin
                        tc = f[625];
                        p[22] = p[22] - tc;
                        p[580] = p[580] + tc;
                end
                627: begin
                        tc = f[626];
                        p[587] = p[587] - tc;
                        p[583] = p[583] + tc;
                end
                628: begin
                        tc = f[627];
                        p[581] = p[581] - tc;
                end
                629: begin
                        tc = f[628];
                        p[585] = p[585] - tc;
                        p[587] = p[587] + tc;
                end
                630: begin
                        tc = f[629];
                        p[582] = p[582] - tc*2;
                        p[588] = p[588] + tc;
                end
                631: begin
                        tc = f[630];
                        p[589] = p[589] - tc;
                        p[586] = p[586] + tc;
                end
                632: begin
                        tc = f[631];
                        p[582] = p[582] - tc;
                        p[591] = p[591] - tc;
                        p[590] = p[590] + tc;
                end
                633: begin
                        tc = f[632];
                        p[592] = p[592] - tc;
                        p[589] = p[589] + tc;
                end
                634: begin
                        tc = f[633];
                        p[581] = p[581] - tc;
                        p[584] = p[584] + tc;
                        p[593] = p[593] + tc;
                end
                635: begin
                        tc = f[634];
                        p[581] = p[581] - tc;
                        p[593] = p[593] + tc;
                end
                636: begin
                        tc = f[635];
                        p[594] = p[594] - tc;
                        p[592] = p[592] + tc;
                end
                637: begin
                        tc = f[636];
                        p[588] = p[588] - tc;
                        p[582] = p[582] + tc;
                end
                638: begin
                        tc = f[637];
                        p[595] = p[595] - tc;
                        p[594] = p[594] + tc;
                end
                639: begin
                        tc = f[638];
                        p[593] = p[593] - tc;
                        p[581] = p[581] + tc*2;
                end
                640: begin
                        tc = f[639];
                        p[583] = p[583] - tc;
                        p[590] = p[590] - tc;
                        p[591] = p[591] + tc;
                        p[595] = p[595] + tc;
                end
                641: begin
                        tc = f[640];
                        p[583] = p[583] - tc;
                        p[595] = p[595] + tc;
                end
                642: begin
                        tc = f[641];
                        p[73] = p[73] - tc;
                        p[581] = p[581] + tc;
                        p[596] = p[596] + tc;
                end
                643: begin
                        tc = f[642];
                        p[596] = p[596] - tc;
                        p[73] = p[73] + tc;
                end
                644: begin
                        tc = f[643];
                        p[598] = p[598] - tc;
                        p[597] = p[597] + tc;
                end
                645: begin
                        tc = f[644];
                        p[599] = p[599] - tc;
                        p[598] = p[598] + tc;
                end
                646: begin
                        tc = f[645];
                        p[74] = p[74] - tc;
                        p[582] = p[582] + tc;
                        p[600] = p[600] + tc;
                end
                647: begin
                        tc = f[646];
                        p[600] = p[600] - tc;
                        p[74] = p[74] + tc;
                end
                648: begin
                        tc = f[647];
                        p[602] = p[602] - tc;
                        p[601] = p[601] + tc;
                end
                649: begin
                        tc = f[648];
                        p[603] = p[603] - tc;
                        p[602] = p[602] + tc;
                end
                650: begin
                        tc = f[649];
                        p[597] = p[597] - tc;
                        p[601] = p[601] - tc;
                        p[22] = p[22] + tc;
                end
                651: begin
                        tc = f[650];
                        p[583] = p[583] - tc;
                        p[599] = p[599] + tc;
                        p[603] = p[603] + tc;
                end
                652: begin
                        tc = f[651];
                        p[584] = p[584] - tc;
                        p[75] = p[75] + tc;
                end
                653: begin
                        tc = f[652];
                        p[75] = p[75] - tc;
                end
                654: begin
                        tc = f[653];
                        p[604] = p[604] - tc;
                        p[585] = p[585] + tc;
                end
                655: begin
                        tc = f[654];
                        p[23] = p[23] - tc;
                        p[604] = p[604] + tc;
                end
                656: begin
                        tc = f[655];
                        p[606] = p[606] - tc;
                        p[607] = p[607] + tc;
                end
                657: begin
                        tc = f[656];
                        p[609] = p[609] - tc;
                        p[608] = p[608] + tc;
                end
                658: begin
                        tc = f[657];
                        p[75] = p[75] - tc;
                        p[605] = p[605] + tc;
                        p[610] = p[610] + tc;
                end
                659: begin
                        tc = f[658];
                        p[610] = p[610] - tc;
                        p[75] = p[75] + tc;
                end
                660: begin
                        tc = f[659];
                        p[612] = p[612] - tc;
                        p[611] = p[611] + tc;
                end
                661: begin
                        tc = f[660];
                        p[613] = p[613] - tc;
                        p[612] = p[612] + tc;
                end
                662: begin
                        tc = f[661];
                        p[70] = p[70] - tc;
                        p[606] = p[606] + tc;
                        p[614] = p[614] + tc;
                end
                663: begin
                        tc = f[662];
                        p[614] = p[614] - tc;
                        p[70] = p[70] + tc;
                end
                664: begin
                        tc = f[663];
                        p[616] = p[616] - tc;
                        p[615] = p[615] + tc;
                end
                665: begin
                        tc = f[664];
                        p[617] = p[617] - tc;
                        p[616] = p[616] + tc;
                end
                666: begin
                        tc = f[665];
                        p[611] = p[611] - tc;
                        p[615] = p[615] - tc;
                        p[23] = p[23] + tc;
                end
                667: begin
                        tc = f[666];
                        p[608] = p[608] - tc;
                        p[613] = p[613] + tc;
                        p[617] = p[617] + tc;
                end
                668: begin
                        tc = f[667];
                        p[607] = p[607] - tc;
                        p[76] = p[76] + tc;
                end
                669: begin
                        tc = f[668];
                        p[76] = p[76] - tc;
                end
                670: begin
                        tc = f[669];
                        p[618] = p[618] - tc;
                        p[609] = p[609] + tc;
                end
                671: begin
                        tc = f[670];
                        p[24] = p[24] - tc;
                        p[618] = p[618] + tc;
                end
                672: begin
                        tc = f[671];
                        p[625] = p[625] - tc;
                        p[621] = p[621] + tc;
                end
                673: begin
                        tc = f[672];
                        p[619] = p[619] - tc;
                end
                674: begin
                        tc = f[673];
                        p[623] = p[623] - tc;
                        p[625] = p[625] + tc;
                end
                675: begin
                        tc = f[674];
                        p[620] = p[620] - tc*2;
                        p[626] = p[626] + tc;
                end
                676: begin
                        tc = f[675];
                        p[627] = p[627] - tc;
                        p[624] = p[624] + tc;
                end
                677: begin
                        tc = f[676];
                        p[620] = p[620] - tc;
                        p[629] = p[629] - tc;
                        p[628] = p[628] + tc;
                end
                678: begin
                        tc = f[677];
                        p[630] = p[630] - tc;
                        p[627] = p[627] + tc;
                end
                679: begin
                        tc = f[678];
                        p[619] = p[619] - tc;
                        p[622] = p[622] + tc;
                        p[631] = p[631] + tc;
                end
                680: begin
                        tc = f[679];
                        p[619] = p[619] - tc;
                        p[631] = p[631] + tc;
                end
                681: begin
                        tc = f[680];
                        p[632] = p[632] - tc;
                        p[630] = p[630] + tc;
                end
                682: begin
                        tc = f[681];
                        p[626] = p[626] - tc;
                        p[620] = p[620] + tc;
                end
                683: begin
                        tc = f[682];
                        p[633] = p[633] - tc;
                        p[632] = p[632] + tc;
                end
                684: begin
                        tc = f[683];
                        p[631] = p[631] - tc;
                        p[619] = p[619] + tc*2;
                end
                685: begin
                        tc = f[684];
                        p[621] = p[621] - tc;
                        p[628] = p[628] - tc;
                        p[629] = p[629] + tc;
                        p[633] = p[633] + tc;
                end
                686: begin
                        tc = f[685];
                        p[621] = p[621] - tc;
                        p[633] = p[633] + tc;
                end
                687: begin
                        tc = f[686];
                        p[77] = p[77] - tc;
                        p[619] = p[619] + tc;
                        p[634] = p[634] + tc;
                end
                688: begin
                        tc = f[687];
                        p[634] = p[634] - tc;
                        p[77] = p[77] + tc;
                end
                689: begin
                        tc = f[688];
                        p[636] = p[636] - tc;
                        p[635] = p[635] + tc;
                end
                690: begin
                        tc = f[689];
                        p[637] = p[637] - tc;
                        p[636] = p[636] + tc;
                end
                691: begin
                        tc = f[690];
                        p[78] = p[78] - tc;
                        p[620] = p[620] + tc;
                        p[638] = p[638] + tc;
                end
                692: begin
                        tc = f[691];
                        p[638] = p[638] - tc;
                        p[78] = p[78] + tc;
                end
                693: begin
                        tc = f[692];
                        p[640] = p[640] - tc;
                        p[639] = p[639] + tc;
                end
                694: begin
                        tc = f[693];
                        p[641] = p[641] - tc;
                        p[640] = p[640] + tc;
                end
                695: begin
                        tc = f[694];
                        p[635] = p[635] - tc;
                        p[639] = p[639] - tc;
                        p[24] = p[24] + tc;
                end
                696: begin
                        tc = f[695];
                        p[621] = p[621] - tc;
                        p[637] = p[637] + tc;
                        p[641] = p[641] + tc;
                end
                697: begin
                        tc = f[696];
                        p[622] = p[622] - tc;
                        p[79] = p[79] + tc;
                end
                698: begin
                        tc = f[697];
                        p[79] = p[79] - tc;
                end
                699: begin
                        tc = f[698];
                        p[642] = p[642] - tc;
                        p[623] = p[623] + tc;
                end
                700: begin
                        tc = f[699];
                        p[25] = p[25] - tc;
                        p[642] = p[642] + tc;
                end
                701: begin
                        tc = f[700];
                        p[644] = p[644] - tc;
                        p[645] = p[645] + tc;
                end
                702: begin
                        tc = f[701];
                        p[647] = p[647] - tc;
                        p[646] = p[646] + tc;
                end
                703: begin
                        tc = f[702];
                        p[79] = p[79] - tc;
                        p[643] = p[643] + tc;
                        p[648] = p[648] + tc;
                end
                704: begin
                        tc = f[703];
                        p[648] = p[648] - tc;
                        p[79] = p[79] + tc;
                end
                705: begin
                        tc = f[704];
                        p[650] = p[650] - tc;
                        p[649] = p[649] + tc;
                end
                706: begin
                        tc = f[705];
                        p[651] = p[651] - tc;
                        p[650] = p[650] + tc;
                end
                707: begin
                        tc = f[706];
                        p[76] = p[76] - tc;
                        p[644] = p[644] + tc;
                        p[652] = p[652] + tc;
                end
                708: begin
                        tc = f[707];
                        p[652] = p[652] - tc;
                        p[76] = p[76] + tc;
                end
                709: begin
                        tc = f[708];
                        p[654] = p[654] - tc;
                        p[653] = p[653] + tc;
                end
                710: begin
                        tc = f[709];
                        p[655] = p[655] - tc;
                        p[654] = p[654] + tc;
                end
                711: begin
                        tc = f[710];
                        p[649] = p[649] - tc;
                        p[653] = p[653] - tc;
                        p[25] = p[25] + tc;
                end
                712: begin
                        tc = f[711];
                        p[646] = p[646] - tc;
                        p[651] = p[651] + tc;
                        p[655] = p[655] + tc;
                end
                713: begin
                        tc = f[712];
                        p[645] = p[645] - tc;
                        p[80] = p[80] + tc;
                end
                714: begin
                        tc = f[713];
                        p[80] = p[80] - tc;
                end
                715: begin
                        tc = f[714];
                        p[656] = p[656] - tc;
                        p[647] = p[647] + tc;
                end
                716: begin
                        tc = f[715];
                        p[26] = p[26] - tc;
                        p[656] = p[656] + tc;
                end
                717: begin
                        tc = f[716];
                        p[658] = p[658] - tc;
                        p[659] = p[659] + tc;
                end
                718: begin
                        tc = f[717];
                        p[661] = p[661] - tc;
                        p[660] = p[660] + tc;
                end
                719: begin
                        tc = f[718];
                        p[80] = p[80] - tc;
                        p[657] = p[657] + tc;
                        p[662] = p[662] + tc;
                end
                720: begin
                        tc = f[719];
                        p[662] = p[662] - tc;
                        p[80] = p[80] + tc;
                end
                721: begin
                        tc = f[720];
                        p[664] = p[664] - tc;
                        p[663] = p[663] + tc;
                end
                722: begin
                        tc = f[721];
                        p[665] = p[665] - tc;
                        p[664] = p[664] + tc;
                end
                723: begin
                        tc = f[722];
                        p[81] = p[81] - tc;
                        p[658] = p[658] + tc;
                        p[666] = p[666] + tc;
                end
                724: begin
                        tc = f[723];
                        p[666] = p[666] - tc;
                        p[81] = p[81] + tc;
                end
                725: begin
                        tc = f[724];
                        p[668] = p[668] - tc;
                        p[667] = p[667] + tc;
                end
                726: begin
                        tc = f[725];
                        p[669] = p[669] - tc;
                        p[668] = p[668] + tc;
                end
                727: begin
                        tc = f[726];
                        p[663] = p[663] - tc;
                        p[667] = p[667] - tc;
                        p[26] = p[26] + tc;
                end
                728: begin
                        tc = f[727];
                        p[660] = p[660] - tc;
                        p[665] = p[665] + tc;
                        p[669] = p[669] + tc;
                end
                729: begin
                        tc = f[728];
                        p[659] = p[659] - tc;
                        p[82] = p[82] + tc;
                end
                730: begin
                        tc = f[729];
                        p[82] = p[82] - tc;
                end
                731: begin
                        tc = f[730];
                        p[670] = p[670] - tc;
                        p[661] = p[661] + tc;
                end
                732: begin
                        tc = f[731];
                        p[27] = p[27] - tc;
                        p[670] = p[670] + tc;
                end
                default:;
        endcase
        led = ~p[82][5:0];
end
endmodule