module sn(
        input clk,
        output reg [5:0] led
);
`define INH(place) ((place) == 0 ? 512 : 0)
reg [9:0] p0=0,p1=1,p2=1,p3=1,p4=1,p5=1,p6=1,p7=1,p8=1,p9=1,p10=1,p11=1,p12=1,p13=1,p14=1,p15=1,p16=1,p17=1,p18=1,p19=1,p20=1,p21=8,p22=2,p23=0,p24=2,p25=0,p26=2,p27=0,p28=2,p29=0,p30=2,p31=0,p32=5,p33=2,p34=0,p35=2,p36=0,p37=2,p38=0,p39=2,p40=0,p41=0,p42=1,p43=2,p44=0,p45=2,p46=0,p47=2,p48=0,p49=0,p50=10,p51=2,p52=0,p53=2,p54=0,p55=0,p56=5,p57=2,p58=0,p59=0,p60=9,p61=0,p62=0,p63=0,p64=1,p65=0,p66=1,p67=1,p68=1,p69=0,p70=1,p71=0,p72=1,p73=1,p74=0,p75=1,p76=1,p77=0,p78=1,p79=1,p80=1,p81=0,p82=1,p83=1,p84=1,p85=1,p86=0,p87=0,p88=1,p89=0,p90=1,p91=1,p92=1,p93=0,p94=1,p95=0,p96=1,p97=1,p98=0,p99=1,p100=1,p101=0,p102=1,p103=1,p104=1,p105=0,p106=1,p107=1,p108=1,p109=1,p110=0,p111=0,p112=1,p113=0,p114=1,p115=1,p116=1,p117=0,p118=1,p119=0,p120=1,p121=1,p122=0,p123=1,p124=1,p125=0,p126=1,p127=1,p128=1,p129=0,p130=1,p131=1,p132=1,p133=1,p134=0,p135=0,p136=1,p137=0,p138=1,p139=1,p140=1,p141=0,p142=1,p143=0,p144=1,p145=1,p146=0,p147=1,p148=1,p149=0,p150=1,p151=1,p152=1,p153=0,p154=1,p155=1,p156=1,p157=1,p158=0,p159=0,p160=1,p161=0,p162=1,p163=1,p164=1,p165=0,p166=1,p167=0,p168=1,p169=1,p170=0,p171=1,p172=1,p173=0,p174=1,p175=1,p176=1,p177=0,p178=1,p179=1,p180=1,p181=1,p182=0,p183=0,p184=1,p185=0,p186=1,p187=1,p188=1,p189=0,p190=1,p191=0,p192=1,p193=1,p194=0,p195=1,p196=1,p197=0,p198=1,p199=1,p200=1,p201=0,p202=1,p203=1,p204=1,p205=1,p206=0,p207=0,p208=1,p209=0,p210=1,p211=1,p212=1,p213=0,p214=1,p215=0,p216=1,p217=1,p218=0,p219=1,p220=1,p221=0,p222=1,p223=1,p224=1,p225=0,p226=1,p227=1,p228=1,p229=1,p230=0,p231=0,p232=1,p233=0,p234=1,p235=1,p236=1,p237=0,p238=1,p239=0,p240=1,p241=1,p242=0,p243=1,p244=1,p245=0,p246=1,p247=1,p248=1,p249=0,p250=1,p251=1,p252=1,p253=1,p254=0,p255=0,p256=1,p257=0,p258=1,p259=1,p260=1,p261=0,p262=1,p263=0,p264=1,p265=1,p266=0,p267=1,p268=1,p269=0,p270=1,p271=1,p272=1,p273=0,p274=1,p275=1,p276=1,p277=1,p278=0,p279=0,p280=0,p281=1,p282=1,p283=0,p284=1,p285=1,p286=1,p287=0,p288=1,p289=1,p290=1,p291=1,p292=0,p293=0,p294=1,p295=0,p296=1,p297=1,p298=1,p299=0,p300=1,p301=0,p302=1,p303=1,p304=0,p305=1,p306=1,p307=0,p308=1,p309=1,p310=1,p311=0,p312=1,p313=1,p314=1,p315=1,p316=0,p317=0,p318=1,p319=0,p320=1,p321=1,p322=1,p323=0,p324=1,p325=0,p326=1,p327=1,p328=0,p329=1,p330=1,p331=0,p332=1,p333=1,p334=1,p335=0,p336=1,p337=1,p338=1,p339=1,p340=0,p341=0,p342=1,p343=0,p344=1,p345=1,p346=1,p347=0,p348=1,p349=0,p350=1,p351=1,p352=0,p353=1,p354=1,p355=0,p356=1,p357=1,p358=1,p359=0,p360=1,p361=1,p362=1,p363=1,p364=0,p365=0,p366=0,p367=1,p368=1,p369=0,p370=1,p371=1,p372=1,p373=0,p374=1,p375=1,p376=1,p377=1,p378=0,p379=0,p380=1,p381=0,p382=1,p383=1,p384=1,p385=0,p386=1,p387=0,p388=1,p389=1,p390=0,p391=1,p392=1,p393=0,p394=1,p395=1,p396=1,p397=0,p398=1,p399=1,p400=1,p401=1,p402=0,p403=0,p404=1,p405=0,p406=1,p407=1,p408=1,p409=0,p410=1,p411=0,p412=1,p413=1,p414=0,p415=1,p416=1,p417=0,p418=1,p419=1,p420=1,p421=0,p422=1,p423=1,p424=1,p425=1,p426=0,p427=0,p428=0,p429=1,p430=1,p431=0,p432=1,p433=1,p434=1,p435=0,p436=1,p437=1,p438=1,p439=1,p440=0,p441=0,p442=1,p443=0,p444=1,p445=1,p446=1,p447=0,p448=1,p449=0,p450=1,p451=1,p452=0,p453=1,p454=1,p455=0,p456=1,p457=1,p458=1,p459=0,p460=1,p461=1,p462=1,p463=1,p464=0,p465=0,p466=0,p467=1,p468=1,p469=0,p470=1,p471=1,p472=1,p473=0,p474=1,p475=1,p476=1,p477=1,p478=0,p479=0,p480=0,p481=1,p482=1,p483=0,p484=1,p485=1,p486=1,p487=0,p488=1,p489=1,p490=1,p491=1;
reg [9:0] f0,f1,f2,f3,f4,f5,f6,f7,f8,f9,f10,f11,f12,f13,f14,f15,f16,f17,f18,f19,f20,f21,f22,f23,f24,f25,f26,f27,f28,f29,f30,f31,f32,f33,f34,f35,f36,f37,f38,f39,f40,f41,f42,f43,f44,f45,f46,f47,f48,f49,f50,f51,f52,f53,f54,f55,f56,f57,f58,f59,f60,f61,f62,f63,f64,f65,f66,f67,f68,f69,f70,f71,f72,f73,f74,f75,f76,f77,f78,f79,f80,f81,f82,f83,f84,f85,f86,f87,f88,f89,f90,f91,f92,f93,f94,f95,f96,f97,f98,f99,f100,f101,f102,f103,f104,f105,f106,f107,f108,f109,f110,f111,f112,f113,f114,f115,f116,f117,f118,f119,f120,f121,f122,f123,f124,f125,f126,f127,f128,f129,f130,f131,f132,f133,f134,f135,f136,f137,f138,f139,f140,f141,f142,f143,f144,f145,f146,f147,f148,f149,f150,f151,f152,f153,f154,f155,f156,f157,f158,f159,f160,f161,f162,f163,f164,f165,f166,f167,f168,f169,f170,f171,f172,f173,f174,f175,f176,f177,f178,f179,f180,f181,f182,f183,f184,f185,f186,f187,f188,f189,f190,f191,f192,f193,f194,f195,f196,f197,f198,f199,f200,f201,f202,f203,f204,f205,f206,f207,f208,f209,f210,f211,f212,f213,f214,f215,f216,f217,f218,f219,f220,f221,f222,f223,f224,f225,f226,f227,f228,f229,f230,f231,f232,f233,f234,f235,f236,f237,f238,f239,f240,f241,f242,f243,f244,f245,f246,f247,f248,f249,f250,f251,f252,f253,f254,f255,f256,f257,f258,f259,f260,f261,f262,f263,f264,f265,f266,f267,f268,f269,f270,f271,f272,f273,f274,f275,f276,f277,f278,f279,f280,f281,f282,f283,f284,f285,f286,f287,f288,f289,f290,f291,f292,f293,f294,f295,f296,f297,f298,f299,f300,f301,f302,f303,f304,f305,f306,f307,f308,f309,f310,f311,f312,f313,f314,f315,f316,f317,f318,f319,f320,f321,f322,f323,f324,f325,f326,f327,f328,f329,f330,f331,f332,f333,f334,f335,f336,f337,f338,f339,f340,f341,f342,f343,f344,f345,f346,f347,f348,f349,f350,f351,f352,f353,f354,f355,f356,f357,f358,f359,f360,f361,f362,f363,f364,f365,f366,f367,f368,f369,f370,f371,f372,f373,f374,f375,f376,f377,f378,f379,f380,f381,f382,f383,f384,f385,f386,f387,f388,f389,f390,f391,f392,f393,f394,f395,f396,f397,f398,f399,f400,f401,f402,f403,f404,f405,f406,f407,f408,f409,f410,f411,f412,f413,f414,f415,f416,f417,f418,f419,f420,f421,f422,f423,f424,f425,f426,f427,f428,f429,f430,f431,f432,f433,f434,f435,f436,f437,f438,f439,f440,f441,f442,f443,f444,f445,f446,f447,f448,f449,f450,f451,f452,f453,f454,f455,f456,f457,f458,f459,f460,f461,f462,f463,f464,f465,f466,f467,f468,f469,f470,f471,f472,f473,f474,f475,f476,f477,f478,f479,f480,f481,f482,f483,f484,f485,f486,f487,f488,f489,f490,f491,f492,f493,f494,f495,f496,f497,f498,f499,f500,f501,f502,f503,f504,f505,f506,f507,f508,f509,f510,f511,f512,f513,f514,f515,f516,f517,f518,f519,f520,f521,f522,f523,f524,f525,f526,f527,f528,f529,f530,f531,f532,f533,f534;
reg [9:0] tf;
reg [9:0] tc;
reg [47:0] counter1=1;
reg [1:0] clk_div; // 2位寄存器用于实现时钟分频

always @(posedge clk) begin
    if(clk_div < 2'b11)
        clk_div <= clk_div + 1; // 计数器自增
    else
        clk_div <= 2'b00; // 重置计数器
end

// 使用clk_div来控制某些逻辑的触发条件
always @(posedge clk) begin
    if (clk_div == 2'b11) begin
        f0 = 512;
        f0 = (f0 >= `INH(p64)) ? `INH(p64) : f0;
        f0 = (f0 > p67) ? p67 : f0;
        f1 = 512;
        f1 = (f1 >= `INH(p88)) ? `INH(p88) : f1;
        f1 = (f1 > p91) ? p91 : f1;
        f2 = 512;
        f2 = (f2 >= `INH(p112)) ? `INH(p112) : f2;
        f2 = (f2 > p115) ? p115 : f2;
        f3 = 512;
        f3 = (f3 >= `INH(p136)) ? `INH(p136) : f3;
        f3 = (f3 > p139) ? p139 : f3;
        f4 = 512;
        f4 = (f4 >= `INH(p160)) ? `INH(p160) : f4;
        f4 = (f4 > p163) ? p163 : f4;
        f5 = 512;
        f5 = (f5 >= `INH(p184)) ? `INH(p184) : f5;
        f5 = (f5 > p187) ? p187 : f5;
        f6 = 512;
        f6 = (f6 >= `INH(p208)) ? `INH(p208) : f6;
        f6 = (f6 > p211) ? p211 : f6;
        f7 = 512;
        f7 = (f7 >= `INH(p232)) ? `INH(p232) : f7;
        f7 = (f7 > p235) ? p235 : f7;
        f8 = 512;
        f8 = (f8 >= `INH(p256)) ? `INH(p256) : f8;
        f8 = (f8 > p259) ? p259 : f8;
        f9 = 512;
        f9 = (f9 > p278) ? p278 : f9;
        f9 = (f9 >= `INH(p281)) ? `INH(p281) : f9;
        f10 = 512;
        f10 = (f10 >= `INH(p294)) ? `INH(p294) : f10;
        f10 = (f10 > p297) ? p297 : f10;
        f11 = 512;
        f11 = (f11 >= `INH(p318)) ? `INH(p318) : f11;
        f11 = (f11 > p321) ? p321 : f11;
        f12 = 512;
        f12 = (f12 >= `INH(p342)) ? `INH(p342) : f12;
        f12 = (f12 > p345) ? p345 : f12;
        f13 = 512;
        f13 = (f13 > p364) ? p364 : f13;
        f13 = (f13 >= `INH(p367)) ? `INH(p367) : f13;
        f14 = 512;
        f14 = (f14 >= `INH(p380)) ? `INH(p380) : f14;
        f14 = (f14 > p383) ? p383 : f14;
        f15 = 512;
        f15 = (f15 >= `INH(p404)) ? `INH(p404) : f15;
        f15 = (f15 > p407) ? p407 : f15;
        f16 = 512;
        f16 = (f16 > p426) ? p426 : f16;
        f16 = (f16 >= `INH(p429)) ? `INH(p429) : f16;
        f17 = 512;
        f17 = (f17 >= `INH(p442)) ? `INH(p442) : f17;
        f17 = (f17 > p445) ? p445 : f17;
        f18 = 512;
        f18 = (f18 > p464) ? p464 : f18;
        f18 = (f18 >= `INH(p467)) ? `INH(p467) : f18;
        f19 = 512;
        f19 = (f19 > p478) ? p478 : f19;
        f19 = (f19 >= `INH(p481)) ? `INH(p481) : f19;
        f20 = 512;
        f20 = (f20 >= `INH(p63)) ? `INH(p63) : f20;
        f20 = (f20 >= `INH(p64)) ? `INH(p64) : f20;
        f20 = (f20 > p68) ? p68 : f20;
        f21 = 512;
        f21 = (f21 > p62) ? p62 : f21;
        f21 = (f21 >= `INH(p68)) ? `INH(p68) : f21;
        f22 = 512;
        f22 = (f22 > p66) ? p66 : f22;
        f22 = (f22 >= `INH(p68)) ? `INH(p68) : f22;
        f23 = 512;
        f23 = (f23 >= p63/2) ? p63/2 : f23;
        f23 = (f23 >= `INH(p67)) ? `INH(p67) : f23;
        f24 = 512;
        f24 = (f24 >= `INH(p67)) ? `INH(p67) : f24;
        f24 = (f24 > p70) ? p70 : f24;
        f25 = 512;
        f25 = (f25 > p63) ? p63 : f25;
        f25 = (f25 >= `INH(p70)) ? `INH(p70) : f25;
        f25 = (f25 > p72) ? p72 : f25;
        f26 = 512;
        f26 = (f26 >= `INH(p70)) ? `INH(p70) : f26;
        f26 = (f26 > p73) ? p73 : f26;
        f27 = 512;
        f27 = (f27 > p62) ? p62 : f27;
        f27 = (f27 >= `INH(p72)) ? `INH(p72) : f27;
        f27 = (f27 >= `INH(p73)) ? `INH(p73) : f27;
        f28 = 512;
        f28 = (f28 > p62) ? p62 : f28;
        f28 = (f28 >= `INH(p71)) ? `INH(p71) : f28;
        f28 = (f28 >= `INH(p73)) ? `INH(p73) : f28;
        f29 = 512;
        f29 = (f29 >= `INH(p73)) ? `INH(p73) : f29;
        f29 = (f29 > p75) ? p75 : f29;
        f30 = 512;
        f30 = (f30 > p69) ? p69 : f30;
        f30 = (f30 >= `INH(p75)) ? `INH(p75) : f30;
        f31 = 512;
        f31 = (f31 >= `INH(p75)) ? `INH(p75) : f31;
        f31 = (f31 > p76) ? p76 : f31;
        f32 = 512;
        f32 = (f32 > p74) ? p74 : f32;
        f32 = (f32 >= `INH(p76)) ? `INH(p76) : f32;
        f33 = 512;
        f33 = (f33 > p64) ? p64 : f33;
        f33 = (f33 > p71) ? p71 : f33;
        f33 = (f33 >= `INH(p72)) ? `INH(p72) : f33;
        f33 = (f33 >= `INH(p76)) ? `INH(p76) : f33;
        f34 = 512;
        f34 = (f34 > p64) ? p64 : f34;
        f34 = (f34 >= `INH(p71)) ? `INH(p71) : f34;
        f34 = (f34 >= `INH(p76)) ? `INH(p76) : f34;
        f35 = 512;
        f35 = (f35 > p21) ? p21 : f35;
        f35 = (f35 >= `INH(p78)) ? `INH(p78) : f35;
        f36 = 512;
        f36 = (f36 > p77) ? p77 : f36;
        f36 = (f36 >= `INH(p79)) ? `INH(p79) : f36;
        f37 = 512;
        f37 = (f37 >= `INH(p21)) ? `INH(p21) : f37;
        f37 = (f37 >= `INH(p78)) ? `INH(p78) : f37;
        f37 = (f37 > p79) ? p79 : f37;
        f38 = 512;
        f38 = (f38 >= `INH(p77)) ? `INH(p77) : f38;
        f38 = (f38 >= `INH(p79)) ? `INH(p79) : f38;
        f38 = (f38 > p80) ? p80 : f38;
        f39 = 512;
        f39 = (f39 > p22) ? p22 : f39;
        f39 = (f39 >= `INH(p82)) ? `INH(p82) : f39;
        f40 = 512;
        f40 = (f40 > p81) ? p81 : f40;
        f40 = (f40 >= `INH(p83)) ? `INH(p83) : f40;
        f41 = 512;
        f41 = (f41 >= `INH(p22)) ? `INH(p22) : f41;
        f41 = (f41 >= `INH(p82)) ? `INH(p82) : f41;
        f41 = (f41 > p83) ? p83 : f41;
        f42 = 512;
        f42 = (f42 >= `INH(p81)) ? `INH(p81) : f42;
        f42 = (f42 >= `INH(p83)) ? `INH(p83) : f42;
        f42 = (f42 > p84) ? p84 : f42;
        f43 = 512;
        f43 = (f43 >= `INH(p0)) ? `INH(p0) : f43;
        f43 = (f43 > p78) ? p78 : f43;
        f43 = (f43 > p82) ? p82 : f43;
        f44 = 512;
        f44 = (f44 > p64) ? p64 : f44;
        f44 = (f44 >= `INH(p80)) ? `INH(p80) : f44;
        f44 = (f44 >= `INH(p84)) ? `INH(p84) : f44;
        f45 = 512;
        f45 = (f45 > p65) ? p65 : f45;
        f45 = (f45 >= `INH(p85)) ? `INH(p85) : f45;
        f46 = 512;
        f46 = (f46 > p23) ? p23 : f46;
        f46 = (f46 >= `INH(p66)) ? `INH(p66) : f46;
        f47 = 512;
        f47 = (f47 >= `INH(p23)) ? `INH(p23) : f47;
        f47 = (f47 >= `INH(p66)) ? `INH(p66) : f47;
        f47 = (f47 > p85) ? p85 : f47;
        f48 = 512;
        f48 = (f48 > p1) ? p1 : f48;
        f48 = (f48 >= `INH(p65)) ? `INH(p65) : f48;
        f48 = (f48 >= `INH(p85)) ? `INH(p85) : f48;
        f49 = 512;
        f49 = (f49 >= `INH(p87)) ? `INH(p87) : f49;
        f49 = (f49 >= `INH(p88)) ? `INH(p88) : f49;
        f49 = (f49 > p92) ? p92 : f49;
        f50 = 512;
        f50 = (f50 > p86) ? p86 : f50;
        f50 = (f50 >= `INH(p92)) ? `INH(p92) : f50;
        f51 = 512;
        f51 = (f51 > p90) ? p90 : f51;
        f51 = (f51 >= `INH(p92)) ? `INH(p92) : f51;
        f52 = 512;
        f52 = (f52 >= p87/2) ? p87/2 : f52;
        f52 = (f52 >= `INH(p91)) ? `INH(p91) : f52;
        f53 = 512;
        f53 = (f53 >= `INH(p91)) ? `INH(p91) : f53;
        f53 = (f53 > p94) ? p94 : f53;
        f54 = 512;
        f54 = (f54 > p87) ? p87 : f54;
        f54 = (f54 >= `INH(p94)) ? `INH(p94) : f54;
        f54 = (f54 > p96) ? p96 : f54;
        f55 = 512;
        f55 = (f55 >= `INH(p94)) ? `INH(p94) : f55;
        f55 = (f55 > p97) ? p97 : f55;
        f56 = 512;
        f56 = (f56 > p86) ? p86 : f56;
        f56 = (f56 >= `INH(p96)) ? `INH(p96) : f56;
        f56 = (f56 >= `INH(p97)) ? `INH(p97) : f56;
        f57 = 512;
        f57 = (f57 > p86) ? p86 : f57;
        f57 = (f57 >= `INH(p95)) ? `INH(p95) : f57;
        f57 = (f57 >= `INH(p97)) ? `INH(p97) : f57;
        f58 = 512;
        f58 = (f58 >= `INH(p97)) ? `INH(p97) : f58;
        f58 = (f58 > p99) ? p99 : f58;
        f59 = 512;
        f59 = (f59 > p93) ? p93 : f59;
        f59 = (f59 >= `INH(p99)) ? `INH(p99) : f59;
        f60 = 512;
        f60 = (f60 >= `INH(p99)) ? `INH(p99) : f60;
        f60 = (f60 > p100) ? p100 : f60;
        f61 = 512;
        f61 = (f61 > p98) ? p98 : f61;
        f61 = (f61 >= `INH(p100)) ? `INH(p100) : f61;
        f62 = 512;
        f62 = (f62 > p88) ? p88 : f62;
        f62 = (f62 > p95) ? p95 : f62;
        f62 = (f62 >= `INH(p96)) ? `INH(p96) : f62;
        f62 = (f62 >= `INH(p100)) ? `INH(p100) : f62;
        f63 = 512;
        f63 = (f63 > p88) ? p88 : f63;
        f63 = (f63 >= `INH(p95)) ? `INH(p95) : f63;
        f63 = (f63 >= `INH(p100)) ? `INH(p100) : f63;
        f64 = 512;
        f64 = (f64 > p23) ? p23 : f64;
        f64 = (f64 >= `INH(p102)) ? `INH(p102) : f64;
        f65 = 512;
        f65 = (f65 > p101) ? p101 : f65;
        f65 = (f65 >= `INH(p103)) ? `INH(p103) : f65;
        f66 = 512;
        f66 = (f66 >= `INH(p23)) ? `INH(p23) : f66;
        f66 = (f66 >= `INH(p102)) ? `INH(p102) : f66;
        f66 = (f66 > p103) ? p103 : f66;
        f67 = 512;
        f67 = (f67 >= `INH(p101)) ? `INH(p101) : f67;
        f67 = (f67 >= `INH(p103)) ? `INH(p103) : f67;
        f67 = (f67 > p104) ? p104 : f67;
        f68 = 512;
        f68 = (f68 > p24) ? p24 : f68;
        f68 = (f68 >= `INH(p106)) ? `INH(p106) : f68;
        f69 = 512;
        f69 = (f69 > p105) ? p105 : f69;
        f69 = (f69 >= `INH(p107)) ? `INH(p107) : f69;
        f70 = 512;
        f70 = (f70 >= `INH(p24)) ? `INH(p24) : f70;
        f70 = (f70 >= `INH(p106)) ? `INH(p106) : f70;
        f70 = (f70 > p107) ? p107 : f70;
        f71 = 512;
        f71 = (f71 >= `INH(p105)) ? `INH(p105) : f71;
        f71 = (f71 >= `INH(p107)) ? `INH(p107) : f71;
        f71 = (f71 > p108) ? p108 : f71;
        f72 = 512;
        f72 = (f72 >= `INH(p1)) ? `INH(p1) : f72;
        f72 = (f72 > p102) ? p102 : f72;
        f72 = (f72 > p106) ? p106 : f72;
        f73 = 512;
        f73 = (f73 > p88) ? p88 : f73;
        f73 = (f73 >= `INH(p104)) ? `INH(p104) : f73;
        f73 = (f73 >= `INH(p108)) ? `INH(p108) : f73;
        f74 = 512;
        f74 = (f74 > p89) ? p89 : f74;
        f74 = (f74 >= `INH(p109)) ? `INH(p109) : f74;
        f75 = 512;
        f75 = (f75 > p25) ? p25 : f75;
        f75 = (f75 >= `INH(p90)) ? `INH(p90) : f75;
        f76 = 512;
        f76 = (f76 >= `INH(p25)) ? `INH(p25) : f76;
        f76 = (f76 >= `INH(p90)) ? `INH(p90) : f76;
        f76 = (f76 > p109) ? p109 : f76;
        f77 = 512;
        f77 = (f77 > p2) ? p2 : f77;
        f77 = (f77 >= `INH(p89)) ? `INH(p89) : f77;
        f77 = (f77 >= `INH(p109)) ? `INH(p109) : f77;
        f78 = 512;
        f78 = (f78 >= `INH(p111)) ? `INH(p111) : f78;
        f78 = (f78 >= `INH(p112)) ? `INH(p112) : f78;
        f78 = (f78 > p116) ? p116 : f78;
        f79 = 512;
        f79 = (f79 > p110) ? p110 : f79;
        f79 = (f79 >= `INH(p116)) ? `INH(p116) : f79;
        f80 = 512;
        f80 = (f80 > p114) ? p114 : f80;
        f80 = (f80 >= `INH(p116)) ? `INH(p116) : f80;
        f81 = 512;
        f81 = (f81 >= p111/2) ? p111/2 : f81;
        f81 = (f81 >= `INH(p115)) ? `INH(p115) : f81;
        f82 = 512;
        f82 = (f82 >= `INH(p115)) ? `INH(p115) : f82;
        f82 = (f82 > p118) ? p118 : f82;
        f83 = 512;
        f83 = (f83 > p111) ? p111 : f83;
        f83 = (f83 >= `INH(p118)) ? `INH(p118) : f83;
        f83 = (f83 > p120) ? p120 : f83;
        f84 = 512;
        f84 = (f84 >= `INH(p118)) ? `INH(p118) : f84;
        f84 = (f84 > p121) ? p121 : f84;
        f85 = 512;
        f85 = (f85 > p110) ? p110 : f85;
        f85 = (f85 >= `INH(p120)) ? `INH(p120) : f85;
        f85 = (f85 >= `INH(p121)) ? `INH(p121) : f85;
        f86 = 512;
        f86 = (f86 > p110) ? p110 : f86;
        f86 = (f86 >= `INH(p119)) ? `INH(p119) : f86;
        f86 = (f86 >= `INH(p121)) ? `INH(p121) : f86;
        f87 = 512;
        f87 = (f87 >= `INH(p121)) ? `INH(p121) : f87;
        f87 = (f87 > p123) ? p123 : f87;
        f88 = 512;
        f88 = (f88 > p117) ? p117 : f88;
        f88 = (f88 >= `INH(p123)) ? `INH(p123) : f88;
        f89 = 512;
        f89 = (f89 >= `INH(p123)) ? `INH(p123) : f89;
        f89 = (f89 > p124) ? p124 : f89;
        f90 = 512;
        f90 = (f90 > p122) ? p122 : f90;
        f90 = (f90 >= `INH(p124)) ? `INH(p124) : f90;
        f91 = 512;
        f91 = (f91 > p112) ? p112 : f91;
        f91 = (f91 > p119) ? p119 : f91;
        f91 = (f91 >= `INH(p120)) ? `INH(p120) : f91;
        f91 = (f91 >= `INH(p124)) ? `INH(p124) : f91;
        f92 = 512;
        f92 = (f92 > p112) ? p112 : f92;
        f92 = (f92 >= `INH(p119)) ? `INH(p119) : f92;
        f92 = (f92 >= `INH(p124)) ? `INH(p124) : f92;
        f93 = 512;
        f93 = (f93 > p25) ? p25 : f93;
        f93 = (f93 >= `INH(p126)) ? `INH(p126) : f93;
        f94 = 512;
        f94 = (f94 > p125) ? p125 : f94;
        f94 = (f94 >= `INH(p127)) ? `INH(p127) : f94;
        f95 = 512;
        f95 = (f95 >= `INH(p25)) ? `INH(p25) : f95;
        f95 = (f95 >= `INH(p126)) ? `INH(p126) : f95;
        f95 = (f95 > p127) ? p127 : f95;
        f96 = 512;
        f96 = (f96 >= `INH(p125)) ? `INH(p125) : f96;
        f96 = (f96 >= `INH(p127)) ? `INH(p127) : f96;
        f96 = (f96 > p128) ? p128 : f96;
        f97 = 512;
        f97 = (f97 > p26) ? p26 : f97;
        f97 = (f97 >= `INH(p130)) ? `INH(p130) : f97;
        f98 = 512;
        f98 = (f98 > p129) ? p129 : f98;
        f98 = (f98 >= `INH(p131)) ? `INH(p131) : f98;
        f99 = 512;
        f99 = (f99 >= `INH(p26)) ? `INH(p26) : f99;
        f99 = (f99 >= `INH(p130)) ? `INH(p130) : f99;
        f99 = (f99 > p131) ? p131 : f99;
        f100 = 512;
        f100 = (f100 >= `INH(p129)) ? `INH(p129) : f100;
        f100 = (f100 >= `INH(p131)) ? `INH(p131) : f100;
        f100 = (f100 > p132) ? p132 : f100;
        f101 = 512;
        f101 = (f101 >= `INH(p2)) ? `INH(p2) : f101;
        f101 = (f101 > p126) ? p126 : f101;
        f101 = (f101 > p130) ? p130 : f101;
        f102 = 512;
        f102 = (f102 > p112) ? p112 : f102;
        f102 = (f102 >= `INH(p128)) ? `INH(p128) : f102;
        f102 = (f102 >= `INH(p132)) ? `INH(p132) : f102;
        f103 = 512;
        f103 = (f103 > p113) ? p113 : f103;
        f103 = (f103 >= `INH(p133)) ? `INH(p133) : f103;
        f104 = 512;
        f104 = (f104 > p27) ? p27 : f104;
        f104 = (f104 >= `INH(p114)) ? `INH(p114) : f104;
        f105 = 512;
        f105 = (f105 >= `INH(p27)) ? `INH(p27) : f105;
        f105 = (f105 >= `INH(p114)) ? `INH(p114) : f105;
        f105 = (f105 > p133) ? p133 : f105;
        f106 = 512;
        f106 = (f106 > p3) ? p3 : f106;
        f106 = (f106 >= `INH(p113)) ? `INH(p113) : f106;
        f106 = (f106 >= `INH(p133)) ? `INH(p133) : f106;
        f107 = 512;
        f107 = (f107 >= `INH(p135)) ? `INH(p135) : f107;
        f107 = (f107 >= `INH(p136)) ? `INH(p136) : f107;
        f107 = (f107 > p140) ? p140 : f107;
        f108 = 512;
        f108 = (f108 > p134) ? p134 : f108;
        f108 = (f108 >= `INH(p140)) ? `INH(p140) : f108;
        f109 = 512;
        f109 = (f109 > p138) ? p138 : f109;
        f109 = (f109 >= `INH(p140)) ? `INH(p140) : f109;
        f110 = 512;
        f110 = (f110 >= p135/2) ? p135/2 : f110;
        f110 = (f110 >= `INH(p139)) ? `INH(p139) : f110;
        f111 = 512;
        f111 = (f111 >= `INH(p139)) ? `INH(p139) : f111;
        f111 = (f111 > p142) ? p142 : f111;
        f112 = 512;
        f112 = (f112 > p135) ? p135 : f112;
        f112 = (f112 >= `INH(p142)) ? `INH(p142) : f112;
        f112 = (f112 > p144) ? p144 : f112;
        f113 = 512;
        f113 = (f113 >= `INH(p142)) ? `INH(p142) : f113;
        f113 = (f113 > p145) ? p145 : f113;
        f114 = 512;
        f114 = (f114 > p134) ? p134 : f114;
        f114 = (f114 >= `INH(p144)) ? `INH(p144) : f114;
        f114 = (f114 >= `INH(p145)) ? `INH(p145) : f114;
        f115 = 512;
        f115 = (f115 > p134) ? p134 : f115;
        f115 = (f115 >= `INH(p143)) ? `INH(p143) : f115;
        f115 = (f115 >= `INH(p145)) ? `INH(p145) : f115;
        f116 = 512;
        f116 = (f116 >= `INH(p145)) ? `INH(p145) : f116;
        f116 = (f116 > p147) ? p147 : f116;
        f117 = 512;
        f117 = (f117 > p141) ? p141 : f117;
        f117 = (f117 >= `INH(p147)) ? `INH(p147) : f117;
        f118 = 512;
        f118 = (f118 >= `INH(p147)) ? `INH(p147) : f118;
        f118 = (f118 > p148) ? p148 : f118;
        f119 = 512;
        f119 = (f119 > p146) ? p146 : f119;
        f119 = (f119 >= `INH(p148)) ? `INH(p148) : f119;
        f120 = 512;
        f120 = (f120 > p136) ? p136 : f120;
        f120 = (f120 > p143) ? p143 : f120;
        f120 = (f120 >= `INH(p144)) ? `INH(p144) : f120;
        f120 = (f120 >= `INH(p148)) ? `INH(p148) : f120;
        f121 = 512;
        f121 = (f121 > p136) ? p136 : f121;
        f121 = (f121 >= `INH(p143)) ? `INH(p143) : f121;
        f121 = (f121 >= `INH(p148)) ? `INH(p148) : f121;
        f122 = 512;
        f122 = (f122 > p27) ? p27 : f122;
        f122 = (f122 >= `INH(p150)) ? `INH(p150) : f122;
        f123 = 512;
        f123 = (f123 > p149) ? p149 : f123;
        f123 = (f123 >= `INH(p151)) ? `INH(p151) : f123;
        f124 = 512;
        f124 = (f124 >= `INH(p27)) ? `INH(p27) : f124;
        f124 = (f124 >= `INH(p150)) ? `INH(p150) : f124;
        f124 = (f124 > p151) ? p151 : f124;
        f125 = 512;
        f125 = (f125 >= `INH(p149)) ? `INH(p149) : f125;
        f125 = (f125 >= `INH(p151)) ? `INH(p151) : f125;
        f125 = (f125 > p152) ? p152 : f125;
        f126 = 512;
        f126 = (f126 > p28) ? p28 : f126;
        f126 = (f126 >= `INH(p154)) ? `INH(p154) : f126;
        f127 = 512;
        f127 = (f127 > p153) ? p153 : f127;
        f127 = (f127 >= `INH(p155)) ? `INH(p155) : f127;
        f128 = 512;
        f128 = (f128 >= `INH(p28)) ? `INH(p28) : f128;
        f128 = (f128 >= `INH(p154)) ? `INH(p154) : f128;
        f128 = (f128 > p155) ? p155 : f128;
        f129 = 512;
        f129 = (f129 >= `INH(p153)) ? `INH(p153) : f129;
        f129 = (f129 >= `INH(p155)) ? `INH(p155) : f129;
        f129 = (f129 > p156) ? p156 : f129;
        f130 = 512;
        f130 = (f130 >= `INH(p3)) ? `INH(p3) : f130;
        f130 = (f130 > p150) ? p150 : f130;
        f130 = (f130 > p154) ? p154 : f130;
        f131 = 512;
        f131 = (f131 > p136) ? p136 : f131;
        f131 = (f131 >= `INH(p152)) ? `INH(p152) : f131;
        f131 = (f131 >= `INH(p156)) ? `INH(p156) : f131;
        f132 = 512;
        f132 = (f132 > p137) ? p137 : f132;
        f132 = (f132 >= `INH(p157)) ? `INH(p157) : f132;
        f133 = 512;
        f133 = (f133 > p29) ? p29 : f133;
        f133 = (f133 >= `INH(p138)) ? `INH(p138) : f133;
        f134 = 512;
        f134 = (f134 >= `INH(p29)) ? `INH(p29) : f134;
        f134 = (f134 >= `INH(p138)) ? `INH(p138) : f134;
        f134 = (f134 > p157) ? p157 : f134;
        f135 = 512;
        f135 = (f135 > p4) ? p4 : f135;
        f135 = (f135 >= `INH(p137)) ? `INH(p137) : f135;
        f135 = (f135 >= `INH(p157)) ? `INH(p157) : f135;
        f136 = 512;
        f136 = (f136 >= `INH(p159)) ? `INH(p159) : f136;
        f136 = (f136 >= `INH(p160)) ? `INH(p160) : f136;
        f136 = (f136 > p164) ? p164 : f136;
        f137 = 512;
        f137 = (f137 > p158) ? p158 : f137;
        f137 = (f137 >= `INH(p164)) ? `INH(p164) : f137;
        f138 = 512;
        f138 = (f138 > p162) ? p162 : f138;
        f138 = (f138 >= `INH(p164)) ? `INH(p164) : f138;
        f139 = 512;
        f139 = (f139 >= p159/2) ? p159/2 : f139;
        f139 = (f139 >= `INH(p163)) ? `INH(p163) : f139;
        f140 = 512;
        f140 = (f140 >= `INH(p163)) ? `INH(p163) : f140;
        f140 = (f140 > p166) ? p166 : f140;
        f141 = 512;
        f141 = (f141 > p159) ? p159 : f141;
        f141 = (f141 >= `INH(p166)) ? `INH(p166) : f141;
        f141 = (f141 > p168) ? p168 : f141;
        f142 = 512;
        f142 = (f142 >= `INH(p166)) ? `INH(p166) : f142;
        f142 = (f142 > p169) ? p169 : f142;
        f143 = 512;
        f143 = (f143 > p158) ? p158 : f143;
        f143 = (f143 >= `INH(p168)) ? `INH(p168) : f143;
        f143 = (f143 >= `INH(p169)) ? `INH(p169) : f143;
        f144 = 512;
        f144 = (f144 > p158) ? p158 : f144;
        f144 = (f144 >= `INH(p167)) ? `INH(p167) : f144;
        f144 = (f144 >= `INH(p169)) ? `INH(p169) : f144;
        f145 = 512;
        f145 = (f145 >= `INH(p169)) ? `INH(p169) : f145;
        f145 = (f145 > p171) ? p171 : f145;
        f146 = 512;
        f146 = (f146 > p165) ? p165 : f146;
        f146 = (f146 >= `INH(p171)) ? `INH(p171) : f146;
        f147 = 512;
        f147 = (f147 >= `INH(p171)) ? `INH(p171) : f147;
        f147 = (f147 > p172) ? p172 : f147;
        f148 = 512;
        f148 = (f148 > p170) ? p170 : f148;
        f148 = (f148 >= `INH(p172)) ? `INH(p172) : f148;
        f149 = 512;
        f149 = (f149 > p160) ? p160 : f149;
        f149 = (f149 > p167) ? p167 : f149;
        f149 = (f149 >= `INH(p168)) ? `INH(p168) : f149;
        f149 = (f149 >= `INH(p172)) ? `INH(p172) : f149;
        f150 = 512;
        f150 = (f150 > p160) ? p160 : f150;
        f150 = (f150 >= `INH(p167)) ? `INH(p167) : f150;
        f150 = (f150 >= `INH(p172)) ? `INH(p172) : f150;
        f151 = 512;
        f151 = (f151 > p29) ? p29 : f151;
        f151 = (f151 >= `INH(p174)) ? `INH(p174) : f151;
        f152 = 512;
        f152 = (f152 > p173) ? p173 : f152;
        f152 = (f152 >= `INH(p175)) ? `INH(p175) : f152;
        f153 = 512;
        f153 = (f153 >= `INH(p29)) ? `INH(p29) : f153;
        f153 = (f153 >= `INH(p174)) ? `INH(p174) : f153;
        f153 = (f153 > p175) ? p175 : f153;
        f154 = 512;
        f154 = (f154 >= `INH(p173)) ? `INH(p173) : f154;
        f154 = (f154 >= `INH(p175)) ? `INH(p175) : f154;
        f154 = (f154 > p176) ? p176 : f154;
        f155 = 512;
        f155 = (f155 > p30) ? p30 : f155;
        f155 = (f155 >= `INH(p178)) ? `INH(p178) : f155;
        f156 = 512;
        f156 = (f156 > p177) ? p177 : f156;
        f156 = (f156 >= `INH(p179)) ? `INH(p179) : f156;
        f157 = 512;
        f157 = (f157 >= `INH(p30)) ? `INH(p30) : f157;
        f157 = (f157 >= `INH(p178)) ? `INH(p178) : f157;
        f157 = (f157 > p179) ? p179 : f157;
        f158 = 512;
        f158 = (f158 >= `INH(p177)) ? `INH(p177) : f158;
        f158 = (f158 >= `INH(p179)) ? `INH(p179) : f158;
        f158 = (f158 > p180) ? p180 : f158;
        f159 = 512;
        f159 = (f159 >= `INH(p4)) ? `INH(p4) : f159;
        f159 = (f159 > p174) ? p174 : f159;
        f159 = (f159 > p178) ? p178 : f159;
        f160 = 512;
        f160 = (f160 > p160) ? p160 : f160;
        f160 = (f160 >= `INH(p176)) ? `INH(p176) : f160;
        f160 = (f160 >= `INH(p180)) ? `INH(p180) : f160;
        f161 = 512;
        f161 = (f161 > p161) ? p161 : f161;
        f161 = (f161 >= `INH(p181)) ? `INH(p181) : f161;
        f162 = 512;
        f162 = (f162 > p31) ? p31 : f162;
        f162 = (f162 >= `INH(p162)) ? `INH(p162) : f162;
        f163 = 512;
        f163 = (f163 >= `INH(p31)) ? `INH(p31) : f163;
        f163 = (f163 >= `INH(p162)) ? `INH(p162) : f163;
        f163 = (f163 > p181) ? p181 : f163;
        f164 = 512;
        f164 = (f164 > p5) ? p5 : f164;
        f164 = (f164 >= `INH(p161)) ? `INH(p161) : f164;
        f164 = (f164 >= `INH(p181)) ? `INH(p181) : f164;
        f165 = 512;
        f165 = (f165 >= `INH(p183)) ? `INH(p183) : f165;
        f165 = (f165 >= `INH(p184)) ? `INH(p184) : f165;
        f165 = (f165 > p188) ? p188 : f165;
        f166 = 512;
        f166 = (f166 > p182) ? p182 : f166;
        f166 = (f166 >= `INH(p188)) ? `INH(p188) : f166;
        f167 = 512;
        f167 = (f167 > p186) ? p186 : f167;
        f167 = (f167 >= `INH(p188)) ? `INH(p188) : f167;
        f168 = 512;
        f168 = (f168 >= p183/2) ? p183/2 : f168;
        f168 = (f168 >= `INH(p187)) ? `INH(p187) : f168;
        f169 = 512;
        f169 = (f169 >= `INH(p187)) ? `INH(p187) : f169;
        f169 = (f169 > p190) ? p190 : f169;
        f170 = 512;
        f170 = (f170 > p183) ? p183 : f170;
        f170 = (f170 >= `INH(p190)) ? `INH(p190) : f170;
        f170 = (f170 > p192) ? p192 : f170;
        f171 = 512;
        f171 = (f171 >= `INH(p190)) ? `INH(p190) : f171;
        f171 = (f171 > p193) ? p193 : f171;
        f172 = 512;
        f172 = (f172 > p182) ? p182 : f172;
        f172 = (f172 >= `INH(p192)) ? `INH(p192) : f172;
        f172 = (f172 >= `INH(p193)) ? `INH(p193) : f172;
        f173 = 512;
        f173 = (f173 > p182) ? p182 : f173;
        f173 = (f173 >= `INH(p191)) ? `INH(p191) : f173;
        f173 = (f173 >= `INH(p193)) ? `INH(p193) : f173;
        f174 = 512;
        f174 = (f174 >= `INH(p193)) ? `INH(p193) : f174;
        f174 = (f174 > p195) ? p195 : f174;
        f175 = 512;
        f175 = (f175 > p189) ? p189 : f175;
        f175 = (f175 >= `INH(p195)) ? `INH(p195) : f175;
        f176 = 512;
        f176 = (f176 >= `INH(p195)) ? `INH(p195) : f176;
        f176 = (f176 > p196) ? p196 : f176;
        f177 = 512;
        f177 = (f177 > p194) ? p194 : f177;
        f177 = (f177 >= `INH(p196)) ? `INH(p196) : f177;
        f178 = 512;
        f178 = (f178 > p184) ? p184 : f178;
        f178 = (f178 > p191) ? p191 : f178;
        f178 = (f178 >= `INH(p192)) ? `INH(p192) : f178;
        f178 = (f178 >= `INH(p196)) ? `INH(p196) : f178;
        f179 = 512;
        f179 = (f179 > p184) ? p184 : f179;
        f179 = (f179 >= `INH(p191)) ? `INH(p191) : f179;
        f179 = (f179 >= `INH(p196)) ? `INH(p196) : f179;
        f180 = 512;
        f180 = (f180 > p32) ? p32 : f180;
        f180 = (f180 >= `INH(p198)) ? `INH(p198) : f180;
        f181 = 512;
        f181 = (f181 > p197) ? p197 : f181;
        f181 = (f181 >= `INH(p199)) ? `INH(p199) : f181;
        f182 = 512;
        f182 = (f182 >= `INH(p32)) ? `INH(p32) : f182;
        f182 = (f182 >= `INH(p198)) ? `INH(p198) : f182;
        f182 = (f182 > p199) ? p199 : f182;
        f183 = 512;
        f183 = (f183 >= `INH(p197)) ? `INH(p197) : f183;
        f183 = (f183 >= `INH(p199)) ? `INH(p199) : f183;
        f183 = (f183 > p200) ? p200 : f183;
        f184 = 512;
        f184 = (f184 > p33) ? p33 : f184;
        f184 = (f184 >= `INH(p202)) ? `INH(p202) : f184;
        f185 = 512;
        f185 = (f185 > p201) ? p201 : f185;
        f185 = (f185 >= `INH(p203)) ? `INH(p203) : f185;
        f186 = 512;
        f186 = (f186 >= `INH(p33)) ? `INH(p33) : f186;
        f186 = (f186 >= `INH(p202)) ? `INH(p202) : f186;
        f186 = (f186 > p203) ? p203 : f186;
        f187 = 512;
        f187 = (f187 >= `INH(p201)) ? `INH(p201) : f187;
        f187 = (f187 >= `INH(p203)) ? `INH(p203) : f187;
        f187 = (f187 > p204) ? p204 : f187;
        f188 = 512;
        f188 = (f188 >= `INH(p5)) ? `INH(p5) : f188;
        f188 = (f188 > p198) ? p198 : f188;
        f188 = (f188 > p202) ? p202 : f188;
        f189 = 512;
        f189 = (f189 > p184) ? p184 : f189;
        f189 = (f189 >= `INH(p200)) ? `INH(p200) : f189;
        f189 = (f189 >= `INH(p204)) ? `INH(p204) : f189;
        f190 = 512;
        f190 = (f190 > p185) ? p185 : f190;
        f190 = (f190 >= `INH(p205)) ? `INH(p205) : f190;
        f191 = 512;
        f191 = (f191 > p34) ? p34 : f191;
        f191 = (f191 >= `INH(p186)) ? `INH(p186) : f191;
        f192 = 512;
        f192 = (f192 >= `INH(p34)) ? `INH(p34) : f192;
        f192 = (f192 >= `INH(p186)) ? `INH(p186) : f192;
        f192 = (f192 > p205) ? p205 : f192;
        f193 = 512;
        f193 = (f193 > p6) ? p6 : f193;
        f193 = (f193 >= `INH(p185)) ? `INH(p185) : f193;
        f193 = (f193 >= `INH(p205)) ? `INH(p205) : f193;
        f194 = 512;
        f194 = (f194 >= `INH(p207)) ? `INH(p207) : f194;
        f194 = (f194 >= `INH(p208)) ? `INH(p208) : f194;
        f194 = (f194 > p212) ? p212 : f194;
        f195 = 512;
        f195 = (f195 > p206) ? p206 : f195;
        f195 = (f195 >= `INH(p212)) ? `INH(p212) : f195;
        f196 = 512;
        f196 = (f196 > p210) ? p210 : f196;
        f196 = (f196 >= `INH(p212)) ? `INH(p212) : f196;
        f197 = 512;
        f197 = (f197 >= p207/2) ? p207/2 : f197;
        f197 = (f197 >= `INH(p211)) ? `INH(p211) : f197;
        f198 = 512;
        f198 = (f198 >= `INH(p211)) ? `INH(p211) : f198;
        f198 = (f198 > p214) ? p214 : f198;
        f199 = 512;
        f199 = (f199 > p207) ? p207 : f199;
        f199 = (f199 >= `INH(p214)) ? `INH(p214) : f199;
        f199 = (f199 > p216) ? p216 : f199;
        f200 = 512;
        f200 = (f200 >= `INH(p214)) ? `INH(p214) : f200;
        f200 = (f200 > p217) ? p217 : f200;
        f201 = 512;
        f201 = (f201 > p206) ? p206 : f201;
        f201 = (f201 >= `INH(p216)) ? `INH(p216) : f201;
        f201 = (f201 >= `INH(p217)) ? `INH(p217) : f201;
        f202 = 512;
        f202 = (f202 > p206) ? p206 : f202;
        f202 = (f202 >= `INH(p215)) ? `INH(p215) : f202;
        f202 = (f202 >= `INH(p217)) ? `INH(p217) : f202;
        f203 = 512;
        f203 = (f203 >= `INH(p217)) ? `INH(p217) : f203;
        f203 = (f203 > p219) ? p219 : f203;
        f204 = 512;
        f204 = (f204 > p213) ? p213 : f204;
        f204 = (f204 >= `INH(p219)) ? `INH(p219) : f204;
        f205 = 512;
        f205 = (f205 >= `INH(p219)) ? `INH(p219) : f205;
        f205 = (f205 > p220) ? p220 : f205;
        f206 = 512;
        f206 = (f206 > p218) ? p218 : f206;
        f206 = (f206 >= `INH(p220)) ? `INH(p220) : f206;
        f207 = 512;
        f207 = (f207 > p208) ? p208 : f207;
        f207 = (f207 > p215) ? p215 : f207;
        f207 = (f207 >= `INH(p216)) ? `INH(p216) : f207;
        f207 = (f207 >= `INH(p220)) ? `INH(p220) : f207;
        f208 = 512;
        f208 = (f208 > p208) ? p208 : f208;
        f208 = (f208 >= `INH(p215)) ? `INH(p215) : f208;
        f208 = (f208 >= `INH(p220)) ? `INH(p220) : f208;
        f209 = 512;
        f209 = (f209 > p34) ? p34 : f209;
        f209 = (f209 >= `INH(p222)) ? `INH(p222) : f209;
        f210 = 512;
        f210 = (f210 > p221) ? p221 : f210;
        f210 = (f210 >= `INH(p223)) ? `INH(p223) : f210;
        f211 = 512;
        f211 = (f211 >= `INH(p34)) ? `INH(p34) : f211;
        f211 = (f211 >= `INH(p222)) ? `INH(p222) : f211;
        f211 = (f211 > p223) ? p223 : f211;
        f212 = 512;
        f212 = (f212 >= `INH(p221)) ? `INH(p221) : f212;
        f212 = (f212 >= `INH(p223)) ? `INH(p223) : f212;
        f212 = (f212 > p224) ? p224 : f212;
        f213 = 512;
        f213 = (f213 > p35) ? p35 : f213;
        f213 = (f213 >= `INH(p226)) ? `INH(p226) : f213;
        f214 = 512;
        f214 = (f214 > p225) ? p225 : f214;
        f214 = (f214 >= `INH(p227)) ? `INH(p227) : f214;
        f215 = 512;
        f215 = (f215 >= `INH(p35)) ? `INH(p35) : f215;
        f215 = (f215 >= `INH(p226)) ? `INH(p226) : f215;
        f215 = (f215 > p227) ? p227 : f215;
        f216 = 512;
        f216 = (f216 >= `INH(p225)) ? `INH(p225) : f216;
        f216 = (f216 >= `INH(p227)) ? `INH(p227) : f216;
        f216 = (f216 > p228) ? p228 : f216;
        f217 = 512;
        f217 = (f217 >= `INH(p6)) ? `INH(p6) : f217;
        f217 = (f217 > p222) ? p222 : f217;
        f217 = (f217 > p226) ? p226 : f217;
        f218 = 512;
        f218 = (f218 > p208) ? p208 : f218;
        f218 = (f218 >= `INH(p224)) ? `INH(p224) : f218;
        f218 = (f218 >= `INH(p228)) ? `INH(p228) : f218;
        f219 = 512;
        f219 = (f219 > p209) ? p209 : f219;
        f219 = (f219 >= `INH(p229)) ? `INH(p229) : f219;
        f220 = 512;
        f220 = (f220 > p36) ? p36 : f220;
        f220 = (f220 >= `INH(p210)) ? `INH(p210) : f220;
        f221 = 512;
        f221 = (f221 >= `INH(p36)) ? `INH(p36) : f221;
        f221 = (f221 >= `INH(p210)) ? `INH(p210) : f221;
        f221 = (f221 > p229) ? p229 : f221;
        f222 = 512;
        f222 = (f222 > p7) ? p7 : f222;
        f222 = (f222 >= `INH(p209)) ? `INH(p209) : f222;
        f222 = (f222 >= `INH(p229)) ? `INH(p229) : f222;
        f223 = 512;
        f223 = (f223 >= `INH(p231)) ? `INH(p231) : f223;
        f223 = (f223 >= `INH(p232)) ? `INH(p232) : f223;
        f223 = (f223 > p236) ? p236 : f223;
        f224 = 512;
        f224 = (f224 > p230) ? p230 : f224;
        f224 = (f224 >= `INH(p236)) ? `INH(p236) : f224;
        f225 = 512;
        f225 = (f225 > p234) ? p234 : f225;
        f225 = (f225 >= `INH(p236)) ? `INH(p236) : f225;
        f226 = 512;
        f226 = (f226 >= p231/2) ? p231/2 : f226;
        f226 = (f226 >= `INH(p235)) ? `INH(p235) : f226;
        f227 = 512;
        f227 = (f227 >= `INH(p235)) ? `INH(p235) : f227;
        f227 = (f227 > p238) ? p238 : f227;
        f228 = 512;
        f228 = (f228 > p231) ? p231 : f228;
        f228 = (f228 >= `INH(p238)) ? `INH(p238) : f228;
        f228 = (f228 > p240) ? p240 : f228;
        f229 = 512;
        f229 = (f229 >= `INH(p238)) ? `INH(p238) : f229;
        f229 = (f229 > p241) ? p241 : f229;
        f230 = 512;
        f230 = (f230 > p230) ? p230 : f230;
        f230 = (f230 >= `INH(p240)) ? `INH(p240) : f230;
        f230 = (f230 >= `INH(p241)) ? `INH(p241) : f230;
        f231 = 512;
        f231 = (f231 > p230) ? p230 : f231;
        f231 = (f231 >= `INH(p239)) ? `INH(p239) : f231;
        f231 = (f231 >= `INH(p241)) ? `INH(p241) : f231;
        f232 = 512;
        f232 = (f232 >= `INH(p241)) ? `INH(p241) : f232;
        f232 = (f232 > p243) ? p243 : f232;
        f233 = 512;
        f233 = (f233 > p237) ? p237 : f233;
        f233 = (f233 >= `INH(p243)) ? `INH(p243) : f233;
        f234 = 512;
        f234 = (f234 >= `INH(p243)) ? `INH(p243) : f234;
        f234 = (f234 > p244) ? p244 : f234;
        f235 = 512;
        f235 = (f235 > p242) ? p242 : f235;
        f235 = (f235 >= `INH(p244)) ? `INH(p244) : f235;
        f236 = 512;
        f236 = (f236 > p232) ? p232 : f236;
        f236 = (f236 > p239) ? p239 : f236;
        f236 = (f236 >= `INH(p240)) ? `INH(p240) : f236;
        f236 = (f236 >= `INH(p244)) ? `INH(p244) : f236;
        f237 = 512;
        f237 = (f237 > p232) ? p232 : f237;
        f237 = (f237 >= `INH(p239)) ? `INH(p239) : f237;
        f237 = (f237 >= `INH(p244)) ? `INH(p244) : f237;
        f238 = 512;
        f238 = (f238 > p36) ? p36 : f238;
        f238 = (f238 >= `INH(p246)) ? `INH(p246) : f238;
        f239 = 512;
        f239 = (f239 > p245) ? p245 : f239;
        f239 = (f239 >= `INH(p247)) ? `INH(p247) : f239;
        f240 = 512;
        f240 = (f240 >= `INH(p36)) ? `INH(p36) : f240;
        f240 = (f240 >= `INH(p246)) ? `INH(p246) : f240;
        f240 = (f240 > p247) ? p247 : f240;
        f241 = 512;
        f241 = (f241 >= `INH(p245)) ? `INH(p245) : f241;
        f241 = (f241 >= `INH(p247)) ? `INH(p247) : f241;
        f241 = (f241 > p248) ? p248 : f241;
        f242 = 512;
        f242 = (f242 > p37) ? p37 : f242;
        f242 = (f242 >= `INH(p250)) ? `INH(p250) : f242;
        f243 = 512;
        f243 = (f243 > p249) ? p249 : f243;
        f243 = (f243 >= `INH(p251)) ? `INH(p251) : f243;
        f244 = 512;
        f244 = (f244 >= `INH(p37)) ? `INH(p37) : f244;
        f244 = (f244 >= `INH(p250)) ? `INH(p250) : f244;
        f244 = (f244 > p251) ? p251 : f244;
        f245 = 512;
        f245 = (f245 >= `INH(p249)) ? `INH(p249) : f245;
        f245 = (f245 >= `INH(p251)) ? `INH(p251) : f245;
        f245 = (f245 > p252) ? p252 : f245;
        f246 = 512;
        f246 = (f246 >= `INH(p7)) ? `INH(p7) : f246;
        f246 = (f246 > p246) ? p246 : f246;
        f246 = (f246 > p250) ? p250 : f246;
        f247 = 512;
        f247 = (f247 > p232) ? p232 : f247;
        f247 = (f247 >= `INH(p248)) ? `INH(p248) : f247;
        f247 = (f247 >= `INH(p252)) ? `INH(p252) : f247;
        f248 = 512;
        f248 = (f248 > p233) ? p233 : f248;
        f248 = (f248 >= `INH(p253)) ? `INH(p253) : f248;
        f249 = 512;
        f249 = (f249 > p38) ? p38 : f249;
        f249 = (f249 >= `INH(p234)) ? `INH(p234) : f249;
        f250 = 512;
        f250 = (f250 >= `INH(p38)) ? `INH(p38) : f250;
        f250 = (f250 >= `INH(p234)) ? `INH(p234) : f250;
        f250 = (f250 > p253) ? p253 : f250;
        f251 = 512;
        f251 = (f251 > p8) ? p8 : f251;
        f251 = (f251 >= `INH(p233)) ? `INH(p233) : f251;
        f251 = (f251 >= `INH(p253)) ? `INH(p253) : f251;
        f252 = 512;
        f252 = (f252 >= `INH(p255)) ? `INH(p255) : f252;
        f252 = (f252 >= `INH(p256)) ? `INH(p256) : f252;
        f252 = (f252 > p260) ? p260 : f252;
        f253 = 512;
        f253 = (f253 > p254) ? p254 : f253;
        f253 = (f253 >= `INH(p260)) ? `INH(p260) : f253;
        f254 = 512;
        f254 = (f254 > p258) ? p258 : f254;
        f254 = (f254 >= `INH(p260)) ? `INH(p260) : f254;
        f255 = 512;
        f255 = (f255 >= p255/2) ? p255/2 : f255;
        f255 = (f255 >= `INH(p259)) ? `INH(p259) : f255;
        f256 = 512;
        f256 = (f256 >= `INH(p259)) ? `INH(p259) : f256;
        f256 = (f256 > p262) ? p262 : f256;
        f257 = 512;
        f257 = (f257 > p255) ? p255 : f257;
        f257 = (f257 >= `INH(p262)) ? `INH(p262) : f257;
        f257 = (f257 > p264) ? p264 : f257;
        f258 = 512;
        f258 = (f258 >= `INH(p262)) ? `INH(p262) : f258;
        f258 = (f258 > p265) ? p265 : f258;
        f259 = 512;
        f259 = (f259 > p254) ? p254 : f259;
        f259 = (f259 >= `INH(p264)) ? `INH(p264) : f259;
        f259 = (f259 >= `INH(p265)) ? `INH(p265) : f259;
        f260 = 512;
        f260 = (f260 > p254) ? p254 : f260;
        f260 = (f260 >= `INH(p263)) ? `INH(p263) : f260;
        f260 = (f260 >= `INH(p265)) ? `INH(p265) : f260;
        f261 = 512;
        f261 = (f261 >= `INH(p265)) ? `INH(p265) : f261;
        f261 = (f261 > p267) ? p267 : f261;
        f262 = 512;
        f262 = (f262 > p261) ? p261 : f262;
        f262 = (f262 >= `INH(p267)) ? `INH(p267) : f262;
        f263 = 512;
        f263 = (f263 >= `INH(p267)) ? `INH(p267) : f263;
        f263 = (f263 > p268) ? p268 : f263;
        f264 = 512;
        f264 = (f264 > p266) ? p266 : f264;
        f264 = (f264 >= `INH(p268)) ? `INH(p268) : f264;
        f265 = 512;
        f265 = (f265 > p256) ? p256 : f265;
        f265 = (f265 > p263) ? p263 : f265;
        f265 = (f265 >= `INH(p264)) ? `INH(p264) : f265;
        f265 = (f265 >= `INH(p268)) ? `INH(p268) : f265;
        f266 = 512;
        f266 = (f266 > p256) ? p256 : f266;
        f266 = (f266 >= `INH(p263)) ? `INH(p263) : f266;
        f266 = (f266 >= `INH(p268)) ? `INH(p268) : f266;
        f267 = 512;
        f267 = (f267 > p38) ? p38 : f267;
        f267 = (f267 >= `INH(p270)) ? `INH(p270) : f267;
        f268 = 512;
        f268 = (f268 > p269) ? p269 : f268;
        f268 = (f268 >= `INH(p271)) ? `INH(p271) : f268;
        f269 = 512;
        f269 = (f269 >= `INH(p38)) ? `INH(p38) : f269;
        f269 = (f269 >= `INH(p270)) ? `INH(p270) : f269;
        f269 = (f269 > p271) ? p271 : f269;
        f270 = 512;
        f270 = (f270 >= `INH(p269)) ? `INH(p269) : f270;
        f270 = (f270 >= `INH(p271)) ? `INH(p271) : f270;
        f270 = (f270 > p272) ? p272 : f270;
        f271 = 512;
        f271 = (f271 > p39) ? p39 : f271;
        f271 = (f271 >= `INH(p274)) ? `INH(p274) : f271;
        f272 = 512;
        f272 = (f272 > p273) ? p273 : f272;
        f272 = (f272 >= `INH(p275)) ? `INH(p275) : f272;
        f273 = 512;
        f273 = (f273 >= `INH(p39)) ? `INH(p39) : f273;
        f273 = (f273 >= `INH(p274)) ? `INH(p274) : f273;
        f273 = (f273 > p275) ? p275 : f273;
        f274 = 512;
        f274 = (f274 >= `INH(p273)) ? `INH(p273) : f274;
        f274 = (f274 >= `INH(p275)) ? `INH(p275) : f274;
        f274 = (f274 > p276) ? p276 : f274;
        f275 = 512;
        f275 = (f275 >= `INH(p8)) ? `INH(p8) : f275;
        f275 = (f275 > p270) ? p270 : f275;
        f275 = (f275 > p274) ? p274 : f275;
        f276 = 512;
        f276 = (f276 > p256) ? p256 : f276;
        f276 = (f276 >= `INH(p272)) ? `INH(p272) : f276;
        f276 = (f276 >= `INH(p276)) ? `INH(p276) : f276;
        f277 = 512;
        f277 = (f277 > p257) ? p257 : f277;
        f277 = (f277 >= `INH(p277)) ? `INH(p277) : f277;
        f278 = 512;
        f278 = (f278 > p40) ? p40 : f278;
        f278 = (f278 >= `INH(p258)) ? `INH(p258) : f278;
        f279 = 512;
        f279 = (f279 >= `INH(p40)) ? `INH(p40) : f279;
        f279 = (f279 >= `INH(p258)) ? `INH(p258) : f279;
        f279 = (f279 > p277) ? p277 : f279;
        f280 = 512;
        f280 = (f280 > p9) ? p9 : f280;
        f280 = (f280 >= `INH(p257)) ? `INH(p257) : f280;
        f280 = (f280 >= `INH(p277)) ? `INH(p277) : f280;
        f281 = 512;
        f281 = (f281 > p279) ? p279 : f281;
        f281 = (f281 >= `INH(p281)) ? `INH(p281) : f281;
        f282 = 512;
        f282 = (f282 >= `INH(p278)) ? `INH(p278) : f282;
        f282 = (f282 >= `INH(p279)) ? `INH(p279) : f282;
        f282 = (f282 >= `INH(p281)) ? `INH(p281) : f282;
        f282 = (f282 > p282) ? p282 : f282;
        f283 = 512;
        f283 = (f283 > p31) ? p31 : f283;
        f283 = (f283 >= `INH(p284)) ? `INH(p284) : f283;
        f284 = 512;
        f284 = (f284 > p283) ? p283 : f284;
        f284 = (f284 >= `INH(p285)) ? `INH(p285) : f284;
        f285 = 512;
        f285 = (f285 >= `INH(p31)) ? `INH(p31) : f285;
        f285 = (f285 >= `INH(p284)) ? `INH(p284) : f285;
        f285 = (f285 > p285) ? p285 : f285;
        f286 = 512;
        f286 = (f286 >= `INH(p283)) ? `INH(p283) : f286;
        f286 = (f286 >= `INH(p285)) ? `INH(p285) : f286;
        f286 = (f286 > p286) ? p286 : f286;
        f287 = 512;
        f287 = (f287 > p40) ? p40 : f287;
        f287 = (f287 >= `INH(p288)) ? `INH(p288) : f287;
        f288 = 512;
        f288 = (f288 > p287) ? p287 : f288;
        f288 = (f288 >= `INH(p289)) ? `INH(p289) : f288;
        f289 = 512;
        f289 = (f289 >= `INH(p40)) ? `INH(p40) : f289;
        f289 = (f289 >= `INH(p288)) ? `INH(p288) : f289;
        f289 = (f289 > p289) ? p289 : f289;
        f290 = 512;
        f290 = (f290 >= `INH(p287)) ? `INH(p287) : f290;
        f290 = (f290 >= `INH(p289)) ? `INH(p289) : f290;
        f290 = (f290 > p290) ? p290 : f290;
        f291 = 512;
        f291 = (f291 >= `INH(p9)) ? `INH(p9) : f291;
        f291 = (f291 > p284) ? p284 : f291;
        f291 = (f291 > p288) ? p288 : f291;
        f292 = 512;
        f292 = (f292 > p281) ? p281 : f292;
        f292 = (f292 >= `INH(p286)) ? `INH(p286) : f292;
        f292 = (f292 >= `INH(p290)) ? `INH(p290) : f292;
        f293 = 512;
        f293 = (f293 > p280) ? p280 : f293;
        f293 = (f293 >= `INH(p291)) ? `INH(p291) : f293;
        f294 = 512;
        f294 = (f294 > p41) ? p41 : f294;
        f294 = (f294 >= `INH(p282)) ? `INH(p282) : f294;
        f295 = 512;
        f295 = (f295 >= `INH(p41)) ? `INH(p41) : f295;
        f295 = (f295 >= `INH(p282)) ? `INH(p282) : f295;
        f295 = (f295 > p291) ? p291 : f295;
        f296 = 512;
        f296 = (f296 > p10) ? p10 : f296;
        f296 = (f296 >= `INH(p280)) ? `INH(p280) : f296;
        f296 = (f296 >= `INH(p291)) ? `INH(p291) : f296;
        f297 = 512;
        f297 = (f297 >= `INH(p293)) ? `INH(p293) : f297;
        f297 = (f297 >= `INH(p294)) ? `INH(p294) : f297;
        f297 = (f297 > p298) ? p298 : f297;
        f298 = 512;
        f298 = (f298 > p292) ? p292 : f298;
        f298 = (f298 >= `INH(p298)) ? `INH(p298) : f298;
        f299 = 512;
        f299 = (f299 > p296) ? p296 : f299;
        f299 = (f299 >= `INH(p298)) ? `INH(p298) : f299;
        f300 = 512;
        f300 = (f300 >= p293/2) ? p293/2 : f300;
        f300 = (f300 >= `INH(p297)) ? `INH(p297) : f300;
        f301 = 512;
        f301 = (f301 >= `INH(p297)) ? `INH(p297) : f301;
        f301 = (f301 > p300) ? p300 : f301;
        f302 = 512;
        f302 = (f302 > p293) ? p293 : f302;
        f302 = (f302 >= `INH(p300)) ? `INH(p300) : f302;
        f302 = (f302 > p302) ? p302 : f302;
        f303 = 512;
        f303 = (f303 >= `INH(p300)) ? `INH(p300) : f303;
        f303 = (f303 > p303) ? p303 : f303;
        f304 = 512;
        f304 = (f304 > p292) ? p292 : f304;
        f304 = (f304 >= `INH(p302)) ? `INH(p302) : f304;
        f304 = (f304 >= `INH(p303)) ? `INH(p303) : f304;
        f305 = 512;
        f305 = (f305 > p292) ? p292 : f305;
        f305 = (f305 >= `INH(p301)) ? `INH(p301) : f305;
        f305 = (f305 >= `INH(p303)) ? `INH(p303) : f305;
        f306 = 512;
        f306 = (f306 >= `INH(p303)) ? `INH(p303) : f306;
        f306 = (f306 > p305) ? p305 : f306;
        f307 = 512;
        f307 = (f307 > p299) ? p299 : f307;
        f307 = (f307 >= `INH(p305)) ? `INH(p305) : f307;
        f308 = 512;
        f308 = (f308 >= `INH(p305)) ? `INH(p305) : f308;
        f308 = (f308 > p306) ? p306 : f308;
        f309 = 512;
        f309 = (f309 > p304) ? p304 : f309;
        f309 = (f309 >= `INH(p306)) ? `INH(p306) : f309;
        f310 = 512;
        f310 = (f310 > p294) ? p294 : f310;
        f310 = (f310 > p301) ? p301 : f310;
        f310 = (f310 >= `INH(p302)) ? `INH(p302) : f310;
        f310 = (f310 >= `INH(p306)) ? `INH(p306) : f310;
        f311 = 512;
        f311 = (f311 > p294) ? p294 : f311;
        f311 = (f311 >= `INH(p301)) ? `INH(p301) : f311;
        f311 = (f311 >= `INH(p306)) ? `INH(p306) : f311;
        f312 = 512;
        f312 = (f312 > p42) ? p42 : f312;
        f312 = (f312 >= `INH(p308)) ? `INH(p308) : f312;
        f313 = 512;
        f313 = (f313 > p307) ? p307 : f313;
        f313 = (f313 >= `INH(p309)) ? `INH(p309) : f313;
        f314 = 512;
        f314 = (f314 >= `INH(p42)) ? `INH(p42) : f314;
        f314 = (f314 >= `INH(p308)) ? `INH(p308) : f314;
        f314 = (f314 > p309) ? p309 : f314;
        f315 = 512;
        f315 = (f315 >= `INH(p307)) ? `INH(p307) : f315;
        f315 = (f315 >= `INH(p309)) ? `INH(p309) : f315;
        f315 = (f315 > p310) ? p310 : f315;
        f316 = 512;
        f316 = (f316 > p43) ? p43 : f316;
        f316 = (f316 >= `INH(p312)) ? `INH(p312) : f316;
        f317 = 512;
        f317 = (f317 > p311) ? p311 : f317;
        f317 = (f317 >= `INH(p313)) ? `INH(p313) : f317;
        f318 = 512;
        f318 = (f318 >= `INH(p43)) ? `INH(p43) : f318;
        f318 = (f318 >= `INH(p312)) ? `INH(p312) : f318;
        f318 = (f318 > p313) ? p313 : f318;
        f319 = 512;
        f319 = (f319 >= `INH(p311)) ? `INH(p311) : f319;
        f319 = (f319 >= `INH(p313)) ? `INH(p313) : f319;
        f319 = (f319 > p314) ? p314 : f319;
        f320 = 512;
        f320 = (f320 >= `INH(p10)) ? `INH(p10) : f320;
        f320 = (f320 > p308) ? p308 : f320;
        f320 = (f320 > p312) ? p312 : f320;
        f321 = 512;
        f321 = (f321 > p294) ? p294 : f321;
        f321 = (f321 >= `INH(p310)) ? `INH(p310) : f321;
        f321 = (f321 >= `INH(p314)) ? `INH(p314) : f321;
        f322 = 512;
        f322 = (f322 > p295) ? p295 : f322;
        f322 = (f322 >= `INH(p315)) ? `INH(p315) : f322;
        f323 = 512;
        f323 = (f323 > p44) ? p44 : f323;
        f323 = (f323 >= `INH(p296)) ? `INH(p296) : f323;
        f324 = 512;
        f324 = (f324 >= `INH(p44)) ? `INH(p44) : f324;
        f324 = (f324 >= `INH(p296)) ? `INH(p296) : f324;
        f324 = (f324 > p315) ? p315 : f324;
        f325 = 512;
        f325 = (f325 > p11) ? p11 : f325;
        f325 = (f325 >= `INH(p295)) ? `INH(p295) : f325;
        f325 = (f325 >= `INH(p315)) ? `INH(p315) : f325;
        f326 = 512;
        f326 = (f326 >= `INH(p317)) ? `INH(p317) : f326;
        f326 = (f326 >= `INH(p318)) ? `INH(p318) : f326;
        f326 = (f326 > p322) ? p322 : f326;
        f327 = 512;
        f327 = (f327 > p316) ? p316 : f327;
        f327 = (f327 >= `INH(p322)) ? `INH(p322) : f327;
        f328 = 512;
        f328 = (f328 > p320) ? p320 : f328;
        f328 = (f328 >= `INH(p322)) ? `INH(p322) : f328;
        f329 = 512;
        f329 = (f329 >= p317/2) ? p317/2 : f329;
        f329 = (f329 >= `INH(p321)) ? `INH(p321) : f329;
        f330 = 512;
        f330 = (f330 >= `INH(p321)) ? `INH(p321) : f330;
        f330 = (f330 > p324) ? p324 : f330;
        f331 = 512;
        f331 = (f331 > p317) ? p317 : f331;
        f331 = (f331 >= `INH(p324)) ? `INH(p324) : f331;
        f331 = (f331 > p326) ? p326 : f331;
        f332 = 512;
        f332 = (f332 >= `INH(p324)) ? `INH(p324) : f332;
        f332 = (f332 > p327) ? p327 : f332;
        f333 = 512;
        f333 = (f333 > p316) ? p316 : f333;
        f333 = (f333 >= `INH(p326)) ? `INH(p326) : f333;
        f333 = (f333 >= `INH(p327)) ? `INH(p327) : f333;
        f334 = 512;
        f334 = (f334 > p316) ? p316 : f334;
        f334 = (f334 >= `INH(p325)) ? `INH(p325) : f334;
        f334 = (f334 >= `INH(p327)) ? `INH(p327) : f334;
        f335 = 512;
        f335 = (f335 >= `INH(p327)) ? `INH(p327) : f335;
        f335 = (f335 > p329) ? p329 : f335;
        f336 = 512;
        f336 = (f336 > p323) ? p323 : f336;
        f336 = (f336 >= `INH(p329)) ? `INH(p329) : f336;
        f337 = 512;
        f337 = (f337 >= `INH(p329)) ? `INH(p329) : f337;
        f337 = (f337 > p330) ? p330 : f337;
        f338 = 512;
        f338 = (f338 > p328) ? p328 : f338;
        f338 = (f338 >= `INH(p330)) ? `INH(p330) : f338;
        f339 = 512;
        f339 = (f339 > p318) ? p318 : f339;
        f339 = (f339 > p325) ? p325 : f339;
        f339 = (f339 >= `INH(p326)) ? `INH(p326) : f339;
        f339 = (f339 >= `INH(p330)) ? `INH(p330) : f339;
        f340 = 512;
        f340 = (f340 > p318) ? p318 : f340;
        f340 = (f340 >= `INH(p325)) ? `INH(p325) : f340;
        f340 = (f340 >= `INH(p330)) ? `INH(p330) : f340;
        f341 = 512;
        f341 = (f341 > p44) ? p44 : f341;
        f341 = (f341 >= `INH(p332)) ? `INH(p332) : f341;
        f342 = 512;
        f342 = (f342 > p331) ? p331 : f342;
        f342 = (f342 >= `INH(p333)) ? `INH(p333) : f342;
        f343 = 512;
        f343 = (f343 >= `INH(p44)) ? `INH(p44) : f343;
        f343 = (f343 >= `INH(p332)) ? `INH(p332) : f343;
        f343 = (f343 > p333) ? p333 : f343;
        f344 = 512;
        f344 = (f344 >= `INH(p331)) ? `INH(p331) : f344;
        f344 = (f344 >= `INH(p333)) ? `INH(p333) : f344;
        f344 = (f344 > p334) ? p334 : f344;
        f345 = 512;
        f345 = (f345 > p45) ? p45 : f345;
        f345 = (f345 >= `INH(p336)) ? `INH(p336) : f345;
        f346 = 512;
        f346 = (f346 > p335) ? p335 : f346;
        f346 = (f346 >= `INH(p337)) ? `INH(p337) : f346;
        f347 = 512;
        f347 = (f347 >= `INH(p45)) ? `INH(p45) : f347;
        f347 = (f347 >= `INH(p336)) ? `INH(p336) : f347;
        f347 = (f347 > p337) ? p337 : f347;
        f348 = 512;
        f348 = (f348 >= `INH(p335)) ? `INH(p335) : f348;
        f348 = (f348 >= `INH(p337)) ? `INH(p337) : f348;
        f348 = (f348 > p338) ? p338 : f348;
        f349 = 512;
        f349 = (f349 >= `INH(p11)) ? `INH(p11) : f349;
        f349 = (f349 > p332) ? p332 : f349;
        f349 = (f349 > p336) ? p336 : f349;
        f350 = 512;
        f350 = (f350 > p318) ? p318 : f350;
        f350 = (f350 >= `INH(p334)) ? `INH(p334) : f350;
        f350 = (f350 >= `INH(p338)) ? `INH(p338) : f350;
        f351 = 512;
        f351 = (f351 > p319) ? p319 : f351;
        f351 = (f351 >= `INH(p339)) ? `INH(p339) : f351;
        f352 = 512;
        f352 = (f352 > p46) ? p46 : f352;
        f352 = (f352 >= `INH(p320)) ? `INH(p320) : f352;
        f353 = 512;
        f353 = (f353 >= `INH(p46)) ? `INH(p46) : f353;
        f353 = (f353 >= `INH(p320)) ? `INH(p320) : f353;
        f353 = (f353 > p339) ? p339 : f353;
        f354 = 512;
        f354 = (f354 > p12) ? p12 : f354;
        f354 = (f354 >= `INH(p319)) ? `INH(p319) : f354;
        f354 = (f354 >= `INH(p339)) ? `INH(p339) : f354;
        f355 = 512;
        f355 = (f355 >= `INH(p341)) ? `INH(p341) : f355;
        f355 = (f355 >= `INH(p342)) ? `INH(p342) : f355;
        f355 = (f355 > p346) ? p346 : f355;
        f356 = 512;
        f356 = (f356 > p340) ? p340 : f356;
        f356 = (f356 >= `INH(p346)) ? `INH(p346) : f356;
        f357 = 512;
        f357 = (f357 > p344) ? p344 : f357;
        f357 = (f357 >= `INH(p346)) ? `INH(p346) : f357;
        f358 = 512;
        f358 = (f358 >= p341/2) ? p341/2 : f358;
        f358 = (f358 >= `INH(p345)) ? `INH(p345) : f358;
        f359 = 512;
        f359 = (f359 >= `INH(p345)) ? `INH(p345) : f359;
        f359 = (f359 > p348) ? p348 : f359;
        f360 = 512;
        f360 = (f360 > p341) ? p341 : f360;
        f360 = (f360 >= `INH(p348)) ? `INH(p348) : f360;
        f360 = (f360 > p350) ? p350 : f360;
        f361 = 512;
        f361 = (f361 >= `INH(p348)) ? `INH(p348) : f361;
        f361 = (f361 > p351) ? p351 : f361;
        f362 = 512;
        f362 = (f362 > p340) ? p340 : f362;
        f362 = (f362 >= `INH(p350)) ? `INH(p350) : f362;
        f362 = (f362 >= `INH(p351)) ? `INH(p351) : f362;
        f363 = 512;
        f363 = (f363 > p340) ? p340 : f363;
        f363 = (f363 >= `INH(p349)) ? `INH(p349) : f363;
        f363 = (f363 >= `INH(p351)) ? `INH(p351) : f363;
        f364 = 512;
        f364 = (f364 >= `INH(p351)) ? `INH(p351) : f364;
        f364 = (f364 > p353) ? p353 : f364;
        f365 = 512;
        f365 = (f365 > p347) ? p347 : f365;
        f365 = (f365 >= `INH(p353)) ? `INH(p353) : f365;
        f366 = 512;
        f366 = (f366 >= `INH(p353)) ? `INH(p353) : f366;
        f366 = (f366 > p354) ? p354 : f366;
        f367 = 512;
        f367 = (f367 > p352) ? p352 : f367;
        f367 = (f367 >= `INH(p354)) ? `INH(p354) : f367;
        f368 = 512;
        f368 = (f368 > p342) ? p342 : f368;
        f368 = (f368 > p349) ? p349 : f368;
        f368 = (f368 >= `INH(p350)) ? `INH(p350) : f368;
        f368 = (f368 >= `INH(p354)) ? `INH(p354) : f368;
        f369 = 512;
        f369 = (f369 > p342) ? p342 : f369;
        f369 = (f369 >= `INH(p349)) ? `INH(p349) : f369;
        f369 = (f369 >= `INH(p354)) ? `INH(p354) : f369;
        f370 = 512;
        f370 = (f370 > p46) ? p46 : f370;
        f370 = (f370 >= `INH(p356)) ? `INH(p356) : f370;
        f371 = 512;
        f371 = (f371 > p355) ? p355 : f371;
        f371 = (f371 >= `INH(p357)) ? `INH(p357) : f371;
        f372 = 512;
        f372 = (f372 >= `INH(p46)) ? `INH(p46) : f372;
        f372 = (f372 >= `INH(p356)) ? `INH(p356) : f372;
        f372 = (f372 > p357) ? p357 : f372;
        f373 = 512;
        f373 = (f373 >= `INH(p355)) ? `INH(p355) : f373;
        f373 = (f373 >= `INH(p357)) ? `INH(p357) : f373;
        f373 = (f373 > p358) ? p358 : f373;
        f374 = 512;
        f374 = (f374 > p47) ? p47 : f374;
        f374 = (f374 >= `INH(p360)) ? `INH(p360) : f374;
        f375 = 512;
        f375 = (f375 > p359) ? p359 : f375;
        f375 = (f375 >= `INH(p361)) ? `INH(p361) : f375;
        f376 = 512;
        f376 = (f376 >= `INH(p47)) ? `INH(p47) : f376;
        f376 = (f376 >= `INH(p360)) ? `INH(p360) : f376;
        f376 = (f376 > p361) ? p361 : f376;
        f377 = 512;
        f377 = (f377 >= `INH(p359)) ? `INH(p359) : f377;
        f377 = (f377 >= `INH(p361)) ? `INH(p361) : f377;
        f377 = (f377 > p362) ? p362 : f377;
        f378 = 512;
        f378 = (f378 >= `INH(p12)) ? `INH(p12) : f378;
        f378 = (f378 > p356) ? p356 : f378;
        f378 = (f378 > p360) ? p360 : f378;
        f379 = 512;
        f379 = (f379 > p342) ? p342 : f379;
        f379 = (f379 >= `INH(p358)) ? `INH(p358) : f379;
        f379 = (f379 >= `INH(p362)) ? `INH(p362) : f379;
        f380 = 512;
        f380 = (f380 > p343) ? p343 : f380;
        f380 = (f380 >= `INH(p363)) ? `INH(p363) : f380;
        f381 = 512;
        f381 = (f381 > p48) ? p48 : f381;
        f381 = (f381 >= `INH(p344)) ? `INH(p344) : f381;
        f382 = 512;
        f382 = (f382 >= `INH(p48)) ? `INH(p48) : f382;
        f382 = (f382 >= `INH(p344)) ? `INH(p344) : f382;
        f382 = (f382 > p363) ? p363 : f382;
        f383 = 512;
        f383 = (f383 > p13) ? p13 : f383;
        f383 = (f383 >= `INH(p343)) ? `INH(p343) : f383;
        f383 = (f383 >= `INH(p363)) ? `INH(p363) : f383;
        f384 = 512;
        f384 = (f384 > p365) ? p365 : f384;
        f384 = (f384 >= `INH(p367)) ? `INH(p367) : f384;
        f385 = 512;
        f385 = (f385 >= `INH(p364)) ? `INH(p364) : f385;
        f385 = (f385 >= `INH(p365)) ? `INH(p365) : f385;
        f385 = (f385 >= `INH(p367)) ? `INH(p367) : f385;
        f385 = (f385 > p368) ? p368 : f385;
        f386 = 512;
        f386 = (f386 > p48) ? p48 : f386;
        f386 = (f386 >= `INH(p370)) ? `INH(p370) : f386;
        f387 = 512;
        f387 = (f387 > p369) ? p369 : f387;
        f387 = (f387 >= `INH(p371)) ? `INH(p371) : f387;
        f388 = 512;
        f388 = (f388 >= `INH(p48)) ? `INH(p48) : f388;
        f388 = (f388 >= `INH(p370)) ? `INH(p370) : f388;
        f388 = (f388 > p371) ? p371 : f388;
        f389 = 512;
        f389 = (f389 >= `INH(p369)) ? `INH(p369) : f389;
        f389 = (f389 >= `INH(p371)) ? `INH(p371) : f389;
        f389 = (f389 > p372) ? p372 : f389;
        f390 = 512;
        f390 = (f390 > p41) ? p41 : f390;
        f390 = (f390 >= `INH(p374)) ? `INH(p374) : f390;
        f391 = 512;
        f391 = (f391 > p373) ? p373 : f391;
        f391 = (f391 >= `INH(p375)) ? `INH(p375) : f391;
        f392 = 512;
        f392 = (f392 >= `INH(p41)) ? `INH(p41) : f392;
        f392 = (f392 >= `INH(p374)) ? `INH(p374) : f392;
        f392 = (f392 > p375) ? p375 : f392;
        f393 = 512;
        f393 = (f393 >= `INH(p373)) ? `INH(p373) : f393;
        f393 = (f393 >= `INH(p375)) ? `INH(p375) : f393;
        f393 = (f393 > p376) ? p376 : f393;
        f394 = 512;
        f394 = (f394 >= `INH(p13)) ? `INH(p13) : f394;
        f394 = (f394 > p370) ? p370 : f394;
        f394 = (f394 > p374) ? p374 : f394;
        f395 = 512;
        f395 = (f395 > p367) ? p367 : f395;
        f395 = (f395 >= `INH(p372)) ? `INH(p372) : f395;
        f395 = (f395 >= `INH(p376)) ? `INH(p376) : f395;
        f396 = 512;
        f396 = (f396 > p366) ? p366 : f396;
        f396 = (f396 >= `INH(p377)) ? `INH(p377) : f396;
        f397 = 512;
        f397 = (f397 > p49) ? p49 : f397;
        f397 = (f397 >= `INH(p368)) ? `INH(p368) : f397;
        f398 = 512;
        f398 = (f398 >= `INH(p49)) ? `INH(p49) : f398;
        f398 = (f398 >= `INH(p368)) ? `INH(p368) : f398;
        f398 = (f398 > p377) ? p377 : f398;
        f399 = 512;
        f399 = (f399 > p14) ? p14 : f399;
        f399 = (f399 >= `INH(p366)) ? `INH(p366) : f399;
        f399 = (f399 >= `INH(p377)) ? `INH(p377) : f399;
        f400 = 512;
        f400 = (f400 >= `INH(p379)) ? `INH(p379) : f400;
        f400 = (f400 >= `INH(p380)) ? `INH(p380) : f400;
        f400 = (f400 > p384) ? p384 : f400;
        f401 = 512;
        f401 = (f401 > p378) ? p378 : f401;
        f401 = (f401 >= `INH(p384)) ? `INH(p384) : f401;
        f402 = 512;
        f402 = (f402 > p382) ? p382 : f402;
        f402 = (f402 >= `INH(p384)) ? `INH(p384) : f402;
        f403 = 512;
        f403 = (f403 >= p379/2) ? p379/2 : f403;
        f403 = (f403 >= `INH(p383)) ? `INH(p383) : f403;
        f404 = 512;
        f404 = (f404 >= `INH(p383)) ? `INH(p383) : f404;
        f404 = (f404 > p386) ? p386 : f404;
        f405 = 512;
        f405 = (f405 > p379) ? p379 : f405;
        f405 = (f405 >= `INH(p386)) ? `INH(p386) : f405;
        f405 = (f405 > p388) ? p388 : f405;
        f406 = 512;
        f406 = (f406 >= `INH(p386)) ? `INH(p386) : f406;
        f406 = (f406 > p389) ? p389 : f406;
        f407 = 512;
        f407 = (f407 > p378) ? p378 : f407;
        f407 = (f407 >= `INH(p388)) ? `INH(p388) : f407;
        f407 = (f407 >= `INH(p389)) ? `INH(p389) : f407;
        f408 = 512;
        f408 = (f408 > p378) ? p378 : f408;
        f408 = (f408 >= `INH(p387)) ? `INH(p387) : f408;
        f408 = (f408 >= `INH(p389)) ? `INH(p389) : f408;
        f409 = 512;
        f409 = (f409 >= `INH(p389)) ? `INH(p389) : f409;
        f409 = (f409 > p391) ? p391 : f409;
        f410 = 512;
        f410 = (f410 > p385) ? p385 : f410;
        f410 = (f410 >= `INH(p391)) ? `INH(p391) : f410;
        f411 = 512;
        f411 = (f411 >= `INH(p391)) ? `INH(p391) : f411;
        f411 = (f411 > p392) ? p392 : f411;
        f412 = 512;
        f412 = (f412 > p390) ? p390 : f412;
        f412 = (f412 >= `INH(p392)) ? `INH(p392) : f412;
        f413 = 512;
        f413 = (f413 > p380) ? p380 : f413;
        f413 = (f413 > p387) ? p387 : f413;
        f413 = (f413 >= `INH(p388)) ? `INH(p388) : f413;
        f413 = (f413 >= `INH(p392)) ? `INH(p392) : f413;
        f414 = 512;
        f414 = (f414 > p380) ? p380 : f414;
        f414 = (f414 >= `INH(p387)) ? `INH(p387) : f414;
        f414 = (f414 >= `INH(p392)) ? `INH(p392) : f414;
        f415 = 512;
        f415 = (f415 > p50) ? p50 : f415;
        f415 = (f415 >= `INH(p394)) ? `INH(p394) : f415;
        f416 = 512;
        f416 = (f416 > p393) ? p393 : f416;
        f416 = (f416 >= `INH(p395)) ? `INH(p395) : f416;
        f417 = 512;
        f417 = (f417 >= `INH(p50)) ? `INH(p50) : f417;
        f417 = (f417 >= `INH(p394)) ? `INH(p394) : f417;
        f417 = (f417 > p395) ? p395 : f417;
        f418 = 512;
        f418 = (f418 >= `INH(p393)) ? `INH(p393) : f418;
        f418 = (f418 >= `INH(p395)) ? `INH(p395) : f418;
        f418 = (f418 > p396) ? p396 : f418;
        f419 = 512;
        f419 = (f419 > p51) ? p51 : f419;
        f419 = (f419 >= `INH(p398)) ? `INH(p398) : f419;
        f420 = 512;
        f420 = (f420 > p397) ? p397 : f420;
        f420 = (f420 >= `INH(p399)) ? `INH(p399) : f420;
        f421 = 512;
        f421 = (f421 >= `INH(p51)) ? `INH(p51) : f421;
        f421 = (f421 >= `INH(p398)) ? `INH(p398) : f421;
        f421 = (f421 > p399) ? p399 : f421;
        f422 = 512;
        f422 = (f422 >= `INH(p397)) ? `INH(p397) : f422;
        f422 = (f422 >= `INH(p399)) ? `INH(p399) : f422;
        f422 = (f422 > p400) ? p400 : f422;
        f423 = 512;
        f423 = (f423 >= `INH(p14)) ? `INH(p14) : f423;
        f423 = (f423 > p394) ? p394 : f423;
        f423 = (f423 > p398) ? p398 : f423;
        f424 = 512;
        f424 = (f424 > p380) ? p380 : f424;
        f424 = (f424 >= `INH(p396)) ? `INH(p396) : f424;
        f424 = (f424 >= `INH(p400)) ? `INH(p400) : f424;
        f425 = 512;
        f425 = (f425 > p381) ? p381 : f425;
        f425 = (f425 >= `INH(p401)) ? `INH(p401) : f425;
        f426 = 512;
        f426 = (f426 > p52) ? p52 : f426;
        f426 = (f426 >= `INH(p382)) ? `INH(p382) : f426;
        f427 = 512;
        f427 = (f427 >= `INH(p52)) ? `INH(p52) : f427;
        f427 = (f427 >= `INH(p382)) ? `INH(p382) : f427;
        f427 = (f427 > p401) ? p401 : f427;
        f428 = 512;
        f428 = (f428 > p15) ? p15 : f428;
        f428 = (f428 >= `INH(p381)) ? `INH(p381) : f428;
        f428 = (f428 >= `INH(p401)) ? `INH(p401) : f428;
        f429 = 512;
        f429 = (f429 >= `INH(p403)) ? `INH(p403) : f429;
        f429 = (f429 >= `INH(p404)) ? `INH(p404) : f429;
        f429 = (f429 > p408) ? p408 : f429;
        f430 = 512;
        f430 = (f430 > p402) ? p402 : f430;
        f430 = (f430 >= `INH(p408)) ? `INH(p408) : f430;
        f431 = 512;
        f431 = (f431 > p406) ? p406 : f431;
        f431 = (f431 >= `INH(p408)) ? `INH(p408) : f431;
        f432 = 512;
        f432 = (f432 >= p403/2) ? p403/2 : f432;
        f432 = (f432 >= `INH(p407)) ? `INH(p407) : f432;
        f433 = 512;
        f433 = (f433 >= `INH(p407)) ? `INH(p407) : f433;
        f433 = (f433 > p410) ? p410 : f433;
        f434 = 512;
        f434 = (f434 > p403) ? p403 : f434;
        f434 = (f434 >= `INH(p410)) ? `INH(p410) : f434;
        f434 = (f434 > p412) ? p412 : f434;
        f435 = 512;
        f435 = (f435 >= `INH(p410)) ? `INH(p410) : f435;
        f435 = (f435 > p413) ? p413 : f435;
        f436 = 512;
        f436 = (f436 > p402) ? p402 : f436;
        f436 = (f436 >= `INH(p412)) ? `INH(p412) : f436;
        f436 = (f436 >= `INH(p413)) ? `INH(p413) : f436;
        f437 = 512;
        f437 = (f437 > p402) ? p402 : f437;
        f437 = (f437 >= `INH(p411)) ? `INH(p411) : f437;
        f437 = (f437 >= `INH(p413)) ? `INH(p413) : f437;
        f438 = 512;
        f438 = (f438 >= `INH(p413)) ? `INH(p413) : f438;
        f438 = (f438 > p415) ? p415 : f438;
        f439 = 512;
        f439 = (f439 > p409) ? p409 : f439;
        f439 = (f439 >= `INH(p415)) ? `INH(p415) : f439;
        f440 = 512;
        f440 = (f440 >= `INH(p415)) ? `INH(p415) : f440;
        f440 = (f440 > p416) ? p416 : f440;
        f441 = 512;
        f441 = (f441 > p414) ? p414 : f441;
        f441 = (f441 >= `INH(p416)) ? `INH(p416) : f441;
        f442 = 512;
        f442 = (f442 > p404) ? p404 : f442;
        f442 = (f442 > p411) ? p411 : f442;
        f442 = (f442 >= `INH(p412)) ? `INH(p412) : f442;
        f442 = (f442 >= `INH(p416)) ? `INH(p416) : f442;
        f443 = 512;
        f443 = (f443 > p404) ? p404 : f443;
        f443 = (f443 >= `INH(p411)) ? `INH(p411) : f443;
        f443 = (f443 >= `INH(p416)) ? `INH(p416) : f443;
        f444 = 512;
        f444 = (f444 > p52) ? p52 : f444;
        f444 = (f444 >= `INH(p418)) ? `INH(p418) : f444;
        f445 = 512;
        f445 = (f445 > p417) ? p417 : f445;
        f445 = (f445 >= `INH(p419)) ? `INH(p419) : f445;
        f446 = 512;
        f446 = (f446 >= `INH(p52)) ? `INH(p52) : f446;
        f446 = (f446 >= `INH(p418)) ? `INH(p418) : f446;
        f446 = (f446 > p419) ? p419 : f446;
        f447 = 512;
        f447 = (f447 >= `INH(p417)) ? `INH(p417) : f447;
        f447 = (f447 >= `INH(p419)) ? `INH(p419) : f447;
        f447 = (f447 > p420) ? p420 : f447;
        f448 = 512;
        f448 = (f448 > p53) ? p53 : f448;
        f448 = (f448 >= `INH(p422)) ? `INH(p422) : f448;
        f449 = 512;
        f449 = (f449 > p421) ? p421 : f449;
        f449 = (f449 >= `INH(p423)) ? `INH(p423) : f449;
        f450 = 512;
        f450 = (f450 >= `INH(p53)) ? `INH(p53) : f450;
        f450 = (f450 >= `INH(p422)) ? `INH(p422) : f450;
        f450 = (f450 > p423) ? p423 : f450;
        f451 = 512;
        f451 = (f451 >= `INH(p421)) ? `INH(p421) : f451;
        f451 = (f451 >= `INH(p423)) ? `INH(p423) : f451;
        f451 = (f451 > p424) ? p424 : f451;
        f452 = 512;
        f452 = (f452 >= `INH(p15)) ? `INH(p15) : f452;
        f452 = (f452 > p418) ? p418 : f452;
        f452 = (f452 > p422) ? p422 : f452;
        f453 = 512;
        f453 = (f453 > p404) ? p404 : f453;
        f453 = (f453 >= `INH(p420)) ? `INH(p420) : f453;
        f453 = (f453 >= `INH(p424)) ? `INH(p424) : f453;
        f454 = 512;
        f454 = (f454 > p405) ? p405 : f454;
        f454 = (f454 >= `INH(p425)) ? `INH(p425) : f454;
        f455 = 512;
        f455 = (f455 > p54) ? p54 : f455;
        f455 = (f455 >= `INH(p406)) ? `INH(p406) : f455;
        f456 = 512;
        f456 = (f456 >= `INH(p54)) ? `INH(p54) : f456;
        f456 = (f456 >= `INH(p406)) ? `INH(p406) : f456;
        f456 = (f456 > p425) ? p425 : f456;
        f457 = 512;
        f457 = (f457 > p16) ? p16 : f457;
        f457 = (f457 >= `INH(p405)) ? `INH(p405) : f457;
        f457 = (f457 >= `INH(p425)) ? `INH(p425) : f457;
        f458 = 512;
        f458 = (f458 > p427) ? p427 : f458;
        f458 = (f458 >= `INH(p429)) ? `INH(p429) : f458;
        f459 = 512;
        f459 = (f459 >= `INH(p426)) ? `INH(p426) : f459;
        f459 = (f459 >= `INH(p427)) ? `INH(p427) : f459;
        f459 = (f459 >= `INH(p429)) ? `INH(p429) : f459;
        f459 = (f459 > p430) ? p430 : f459;
        f460 = 512;
        f460 = (f460 > p54) ? p54 : f460;
        f460 = (f460 >= `INH(p432)) ? `INH(p432) : f460;
        f461 = 512;
        f461 = (f461 > p431) ? p431 : f461;
        f461 = (f461 >= `INH(p433)) ? `INH(p433) : f461;
        f462 = 512;
        f462 = (f462 >= `INH(p54)) ? `INH(p54) : f462;
        f462 = (f462 >= `INH(p432)) ? `INH(p432) : f462;
        f462 = (f462 > p433) ? p433 : f462;
        f463 = 512;
        f463 = (f463 >= `INH(p431)) ? `INH(p431) : f463;
        f463 = (f463 >= `INH(p433)) ? `INH(p433) : f463;
        f463 = (f463 > p434) ? p434 : f463;
        f464 = 512;
        f464 = (f464 > p49) ? p49 : f464;
        f464 = (f464 >= `INH(p436)) ? `INH(p436) : f464;
        f465 = 512;
        f465 = (f465 > p435) ? p435 : f465;
        f465 = (f465 >= `INH(p437)) ? `INH(p437) : f465;
        f466 = 512;
        f466 = (f466 >= `INH(p49)) ? `INH(p49) : f466;
        f466 = (f466 >= `INH(p436)) ? `INH(p436) : f466;
        f466 = (f466 > p437) ? p437 : f466;
        f467 = 512;
        f467 = (f467 >= `INH(p435)) ? `INH(p435) : f467;
        f467 = (f467 >= `INH(p437)) ? `INH(p437) : f467;
        f467 = (f467 > p438) ? p438 : f467;
        f468 = 512;
        f468 = (f468 >= `INH(p16)) ? `INH(p16) : f468;
        f468 = (f468 > p432) ? p432 : f468;
        f468 = (f468 > p436) ? p436 : f468;
        f469 = 512;
        f469 = (f469 > p429) ? p429 : f469;
        f469 = (f469 >= `INH(p434)) ? `INH(p434) : f469;
        f469 = (f469 >= `INH(p438)) ? `INH(p438) : f469;
        f470 = 512;
        f470 = (f470 > p428) ? p428 : f470;
        f470 = (f470 >= `INH(p439)) ? `INH(p439) : f470;
        f471 = 512;
        f471 = (f471 > p55) ? p55 : f471;
        f471 = (f471 >= `INH(p430)) ? `INH(p430) : f471;
        f472 = 512;
        f472 = (f472 >= `INH(p55)) ? `INH(p55) : f472;
        f472 = (f472 >= `INH(p430)) ? `INH(p430) : f472;
        f472 = (f472 > p439) ? p439 : f472;
        f473 = 512;
        f473 = (f473 > p17) ? p17 : f473;
        f473 = (f473 >= `INH(p428)) ? `INH(p428) : f473;
        f473 = (f473 >= `INH(p439)) ? `INH(p439) : f473;
        f474 = 512;
        f474 = (f474 >= `INH(p441)) ? `INH(p441) : f474;
        f474 = (f474 >= `INH(p442)) ? `INH(p442) : f474;
        f474 = (f474 > p446) ? p446 : f474;
        f475 = 512;
        f475 = (f475 > p440) ? p440 : f475;
        f475 = (f475 >= `INH(p446)) ? `INH(p446) : f475;
        f476 = 512;
        f476 = (f476 > p444) ? p444 : f476;
        f476 = (f476 >= `INH(p446)) ? `INH(p446) : f476;
        f477 = 512;
        f477 = (f477 >= p441/2) ? p441/2 : f477;
        f477 = (f477 >= `INH(p445)) ? `INH(p445) : f477;
        f478 = 512;
        f478 = (f478 >= `INH(p445)) ? `INH(p445) : f478;
        f478 = (f478 > p448) ? p448 : f478;
        f479 = 512;
        f479 = (f479 > p441) ? p441 : f479;
        f479 = (f479 >= `INH(p448)) ? `INH(p448) : f479;
        f479 = (f479 > p450) ? p450 : f479;
        f480 = 512;
        f480 = (f480 >= `INH(p448)) ? `INH(p448) : f480;
        f480 = (f480 > p451) ? p451 : f480;
        f481 = 512;
        f481 = (f481 > p440) ? p440 : f481;
        f481 = (f481 >= `INH(p450)) ? `INH(p450) : f481;
        f481 = (f481 >= `INH(p451)) ? `INH(p451) : f481;
        f482 = 512;
        f482 = (f482 > p440) ? p440 : f482;
        f482 = (f482 >= `INH(p449)) ? `INH(p449) : f482;
        f482 = (f482 >= `INH(p451)) ? `INH(p451) : f482;
        f483 = 512;
        f483 = (f483 >= `INH(p451)) ? `INH(p451) : f483;
        f483 = (f483 > p453) ? p453 : f483;
        f484 = 512;
        f484 = (f484 > p447) ? p447 : f484;
        f484 = (f484 >= `INH(p453)) ? `INH(p453) : f484;
        f485 = 512;
        f485 = (f485 >= `INH(p453)) ? `INH(p453) : f485;
        f485 = (f485 > p454) ? p454 : f485;
        f486 = 512;
        f486 = (f486 > p452) ? p452 : f486;
        f486 = (f486 >= `INH(p454)) ? `INH(p454) : f486;
        f487 = 512;
        f487 = (f487 > p442) ? p442 : f487;
        f487 = (f487 > p449) ? p449 : f487;
        f487 = (f487 >= `INH(p450)) ? `INH(p450) : f487;
        f487 = (f487 >= `INH(p454)) ? `INH(p454) : f487;
        f488 = 512;
        f488 = (f488 > p442) ? p442 : f488;
        f488 = (f488 >= `INH(p449)) ? `INH(p449) : f488;
        f488 = (f488 >= `INH(p454)) ? `INH(p454) : f488;
        f489 = 512;
        f489 = (f489 > p56) ? p56 : f489;
        f489 = (f489 >= `INH(p456)) ? `INH(p456) : f489;
        f490 = 512;
        f490 = (f490 > p455) ? p455 : f490;
        f490 = (f490 >= `INH(p457)) ? `INH(p457) : f490;
        f491 = 512;
        f491 = (f491 >= `INH(p56)) ? `INH(p56) : f491;
        f491 = (f491 >= `INH(p456)) ? `INH(p456) : f491;
        f491 = (f491 > p457) ? p457 : f491;
        f492 = 512;
        f492 = (f492 >= `INH(p455)) ? `INH(p455) : f492;
        f492 = (f492 >= `INH(p457)) ? `INH(p457) : f492;
        f492 = (f492 > p458) ? p458 : f492;
        f493 = 512;
        f493 = (f493 > p57) ? p57 : f493;
        f493 = (f493 >= `INH(p460)) ? `INH(p460) : f493;
        f494 = 512;
        f494 = (f494 > p459) ? p459 : f494;
        f494 = (f494 >= `INH(p461)) ? `INH(p461) : f494;
        f495 = 512;
        f495 = (f495 >= `INH(p57)) ? `INH(p57) : f495;
        f495 = (f495 >= `INH(p460)) ? `INH(p460) : f495;
        f495 = (f495 > p461) ? p461 : f495;
        f496 = 512;
        f496 = (f496 >= `INH(p459)) ? `INH(p459) : f496;
        f496 = (f496 >= `INH(p461)) ? `INH(p461) : f496;
        f496 = (f496 > p462) ? p462 : f496;
        f497 = 512;
        f497 = (f497 >= `INH(p17)) ? `INH(p17) : f497;
        f497 = (f497 > p456) ? p456 : f497;
        f497 = (f497 > p460) ? p460 : f497;
        f498 = 512;
        f498 = (f498 > p442) ? p442 : f498;
        f498 = (f498 >= `INH(p458)) ? `INH(p458) : f498;
        f498 = (f498 >= `INH(p462)) ? `INH(p462) : f498;
        f499 = 512;
        f499 = (f499 > p443) ? p443 : f499;
        f499 = (f499 >= `INH(p463)) ? `INH(p463) : f499;
        f500 = 512;
        f500 = (f500 > p58) ? p58 : f500;
        f500 = (f500 >= `INH(p444)) ? `INH(p444) : f500;
        f501 = 512;
        f501 = (f501 >= `INH(p58)) ? `INH(p58) : f501;
        f501 = (f501 >= `INH(p444)) ? `INH(p444) : f501;
        f501 = (f501 > p463) ? p463 : f501;
        f502 = 512;
        f502 = (f502 > p18) ? p18 : f502;
        f502 = (f502 >= `INH(p443)) ? `INH(p443) : f502;
        f502 = (f502 >= `INH(p463)) ? `INH(p463) : f502;
        f503 = 512;
        f503 = (f503 > p465) ? p465 : f503;
        f503 = (f503 >= `INH(p467)) ? `INH(p467) : f503;
        f504 = 512;
        f504 = (f504 >= `INH(p464)) ? `INH(p464) : f504;
        f504 = (f504 >= `INH(p465)) ? `INH(p465) : f504;
        f504 = (f504 >= `INH(p467)) ? `INH(p467) : f504;
        f504 = (f504 > p468) ? p468 : f504;
        f505 = 512;
        f505 = (f505 > p58) ? p58 : f505;
        f505 = (f505 >= `INH(p470)) ? `INH(p470) : f505;
        f506 = 512;
        f506 = (f506 > p469) ? p469 : f506;
        f506 = (f506 >= `INH(p471)) ? `INH(p471) : f506;
        f507 = 512;
        f507 = (f507 >= `INH(p58)) ? `INH(p58) : f507;
        f507 = (f507 >= `INH(p470)) ? `INH(p470) : f507;
        f507 = (f507 > p471) ? p471 : f507;
        f508 = 512;
        f508 = (f508 >= `INH(p469)) ? `INH(p469) : f508;
        f508 = (f508 >= `INH(p471)) ? `INH(p471) : f508;
        f508 = (f508 > p472) ? p472 : f508;
        f509 = 512;
        f509 = (f509 > p55) ? p55 : f509;
        f509 = (f509 >= `INH(p474)) ? `INH(p474) : f509;
        f510 = 512;
        f510 = (f510 > p473) ? p473 : f510;
        f510 = (f510 >= `INH(p475)) ? `INH(p475) : f510;
        f511 = 512;
        f511 = (f511 >= `INH(p55)) ? `INH(p55) : f511;
        f511 = (f511 >= `INH(p474)) ? `INH(p474) : f511;
        f511 = (f511 > p475) ? p475 : f511;
        f512 = 512;
        f512 = (f512 >= `INH(p473)) ? `INH(p473) : f512;
        f512 = (f512 >= `INH(p475)) ? `INH(p475) : f512;
        f512 = (f512 > p476) ? p476 : f512;
        f513 = 512;
        f513 = (f513 >= `INH(p18)) ? `INH(p18) : f513;
        f513 = (f513 > p470) ? p470 : f513;
        f513 = (f513 > p474) ? p474 : f513;
        f514 = 512;
        f514 = (f514 > p467) ? p467 : f514;
        f514 = (f514 >= `INH(p472)) ? `INH(p472) : f514;
        f514 = (f514 >= `INH(p476)) ? `INH(p476) : f514;
        f515 = 512;
        f515 = (f515 > p466) ? p466 : f515;
        f515 = (f515 >= `INH(p477)) ? `INH(p477) : f515;
        f516 = 512;
        f516 = (f516 > p59) ? p59 : f516;
        f516 = (f516 >= `INH(p468)) ? `INH(p468) : f516;
        f517 = 512;
        f517 = (f517 >= `INH(p59)) ? `INH(p59) : f517;
        f517 = (f517 >= `INH(p468)) ? `INH(p468) : f517;
        f517 = (f517 > p477) ? p477 : f517;
        f518 = 512;
        f518 = (f518 > p19) ? p19 : f518;
        f518 = (f518 >= `INH(p466)) ? `INH(p466) : f518;
        f518 = (f518 >= `INH(p477)) ? `INH(p477) : f518;
        f519 = 512;
        f519 = (f519 > p479) ? p479 : f519;
        f519 = (f519 >= `INH(p481)) ? `INH(p481) : f519;
        f520 = 512;
        f520 = (f520 >= `INH(p478)) ? `INH(p478) : f520;
        f520 = (f520 >= `INH(p479)) ? `INH(p479) : f520;
        f520 = (f520 >= `INH(p481)) ? `INH(p481) : f520;
        f520 = (f520 > p482) ? p482 : f520;
        f521 = 512;
        f521 = (f521 > p59) ? p59 : f521;
        f521 = (f521 >= `INH(p484)) ? `INH(p484) : f521;
        f522 = 512;
        f522 = (f522 > p483) ? p483 : f522;
        f522 = (f522 >= `INH(p485)) ? `INH(p485) : f522;
        f523 = 512;
        f523 = (f523 >= `INH(p59)) ? `INH(p59) : f523;
        f523 = (f523 >= `INH(p484)) ? `INH(p484) : f523;
        f523 = (f523 > p485) ? p485 : f523;
        f524 = 512;
        f524 = (f524 >= `INH(p483)) ? `INH(p483) : f524;
        f524 = (f524 >= `INH(p485)) ? `INH(p485) : f524;
        f524 = (f524 > p486) ? p486 : f524;
        f525 = 512;
        f525 = (f525 > p60) ? p60 : f525;
        f525 = (f525 >= `INH(p488)) ? `INH(p488) : f525;
        f526 = 512;
        f526 = (f526 > p487) ? p487 : f526;
        f526 = (f526 >= `INH(p489)) ? `INH(p489) : f526;
        f527 = 512;
        f527 = (f527 >= `INH(p60)) ? `INH(p60) : f527;
        f527 = (f527 >= `INH(p488)) ? `INH(p488) : f527;
        f527 = (f527 > p489) ? p489 : f527;
        f528 = 512;
        f528 = (f528 >= `INH(p487)) ? `INH(p487) : f528;
        f528 = (f528 >= `INH(p489)) ? `INH(p489) : f528;
        f528 = (f528 > p490) ? p490 : f528;
        f529 = 512;
        f529 = (f529 >= `INH(p19)) ? `INH(p19) : f529;
        f529 = (f529 > p484) ? p484 : f529;
        f529 = (f529 > p488) ? p488 : f529;
        f530 = 512;
        f530 = (f530 > p481) ? p481 : f530;
        f530 = (f530 >= `INH(p486)) ? `INH(p486) : f530;
        f530 = (f530 >= `INH(p490)) ? `INH(p490) : f530;
        f531 = 512;
        f531 = (f531 > p480) ? p480 : f531;
        f531 = (f531 >= `INH(p491)) ? `INH(p491) : f531;
        f532 = 512;
        f532 = (f532 > p61) ? p61 : f532;
        f532 = (f532 >= `INH(p482)) ? `INH(p482) : f532;
        f533 = 512;
        f533 = (f533 >= `INH(p61)) ? `INH(p61) : f533;
        f533 = (f533 >= `INH(p482)) ? `INH(p482) : f533;
        f533 = (f533 > p491) ? p491 : f533;
        f534 = 512;
        f534 = (f534 > p20) ? p20 : f534;
        f534 = (f534 >= `INH(p480)) ? `INH(p480) : f534;
        f534 = (f534 >= `INH(p491)) ? `INH(p491) : f534;
        if(f20>0)
                f0 = 0;
        if(f21>0)
                f22 = 0;
        if(f23>0)
                f24 = 0;
        if(f25>0)
                f26 = 0;
        if(f27>0)
                f29 = 0;
        if(f28>0)
                f29 = 0;
        if(f30>0)
                f31 = 0;
        if(f32>0)
                f33 = 0;
        if(f32>0)
                f34 = 0;
        if(f49>0)
                f1 = 0;
        if(f50>0)
                f51 = 0;
        if(f52>0)
                f53 = 0;
        if(f54>0)
                f55 = 0;
        if(f56>0)
                f58 = 0;
        if(f57>0)
                f58 = 0;
        if(f59>0)
                f60 = 0;
        if(f61>0)
                f62 = 0;
        if(f61>0)
                f63 = 0;
        if(f78>0)
                f2 = 0;
        if(f79>0)
                f80 = 0;
        if(f81>0)
                f82 = 0;
        if(f83>0)
                f84 = 0;
        if(f85>0)
                f87 = 0;
        if(f86>0)
                f87 = 0;
        if(f88>0)
                f89 = 0;
        if(f90>0)
                f91 = 0;
        if(f90>0)
                f92 = 0;
        if(f107>0)
                f3 = 0;
        if(f108>0)
                f109 = 0;
        if(f110>0)
                f111 = 0;
        if(f112>0)
                f113 = 0;
        if(f114>0)
                f116 = 0;
        if(f115>0)
                f116 = 0;
        if(f117>0)
                f118 = 0;
        if(f119>0)
                f120 = 0;
        if(f119>0)
                f121 = 0;
        if(f136>0)
                f4 = 0;
        if(f137>0)
                f138 = 0;
        if(f139>0)
                f140 = 0;
        if(f141>0)
                f142 = 0;
        if(f143>0)
                f145 = 0;
        if(f144>0)
                f145 = 0;
        if(f146>0)
                f147 = 0;
        if(f148>0)
                f149 = 0;
        if(f148>0)
                f150 = 0;
        if(f165>0)
                f5 = 0;
        if(f166>0)
                f167 = 0;
        if(f168>0)
                f169 = 0;
        if(f170>0)
                f171 = 0;
        if(f172>0)
                f174 = 0;
        if(f173>0)
                f174 = 0;
        if(f175>0)
                f176 = 0;
        if(f177>0)
                f178 = 0;
        if(f177>0)
                f179 = 0;
        if(f194>0)
                f6 = 0;
        if(f195>0)
                f196 = 0;
        if(f197>0)
                f198 = 0;
        if(f199>0)
                f200 = 0;
        if(f201>0)
                f203 = 0;
        if(f202>0)
                f203 = 0;
        if(f204>0)
                f205 = 0;
        if(f206>0)
                f207 = 0;
        if(f206>0)
                f208 = 0;
        if(f223>0)
                f7 = 0;
        if(f224>0)
                f225 = 0;
        if(f226>0)
                f227 = 0;
        if(f228>0)
                f229 = 0;
        if(f230>0)
                f232 = 0;
        if(f231>0)
                f232 = 0;
        if(f233>0)
                f234 = 0;
        if(f235>0)
                f236 = 0;
        if(f235>0)
                f237 = 0;
        if(f252>0)
                f8 = 0;
        if(f253>0)
                f254 = 0;
        if(f255>0)
                f256 = 0;
        if(f257>0)
                f258 = 0;
        if(f259>0)
                f261 = 0;
        if(f260>0)
                f261 = 0;
        if(f262>0)
                f263 = 0;
        if(f264>0)
                f265 = 0;
        if(f264>0)
                f266 = 0;
        if(f297>0)
                f10 = 0;
        if(f298>0)
                f299 = 0;
        if(f300>0)
                f301 = 0;
        if(f302>0)
                f303 = 0;
        if(f304>0)
                f306 = 0;
        if(f305>0)
                f306 = 0;
        if(f307>0)
                f308 = 0;
        if(f309>0)
                f310 = 0;
        if(f309>0)
                f311 = 0;
        if(f326>0)
                f11 = 0;
        if(f327>0)
                f328 = 0;
        if(f329>0)
                f330 = 0;
        if(f331>0)
                f332 = 0;
        if(f333>0)
                f335 = 0;
        if(f334>0)
                f335 = 0;
        if(f336>0)
                f337 = 0;
        if(f338>0)
                f339 = 0;
        if(f338>0)
                f340 = 0;
        if(f355>0)
                f12 = 0;
        if(f356>0)
                f357 = 0;
        if(f358>0)
                f359 = 0;
        if(f360>0)
                f361 = 0;
        if(f362>0)
                f364 = 0;
        if(f363>0)
                f364 = 0;
        if(f365>0)
                f366 = 0;
        if(f367>0)
                f368 = 0;
        if(f367>0)
                f369 = 0;
        if(f400>0)
                f14 = 0;
        if(f401>0)
                f402 = 0;
        if(f403>0)
                f404 = 0;
        if(f405>0)
                f406 = 0;
        if(f407>0)
                f409 = 0;
        if(f408>0)
                f409 = 0;
        if(f410>0)
                f411 = 0;
        if(f412>0)
                f413 = 0;
        if(f412>0)
                f414 = 0;
        if(f429>0)
                f15 = 0;
        if(f430>0)
                f431 = 0;
        if(f432>0)
                f433 = 0;
        if(f434>0)
                f435 = 0;
        if(f436>0)
                f438 = 0;
        if(f437>0)
                f438 = 0;
        if(f439>0)
                f440 = 0;
        if(f441>0)
                f442 = 0;
        if(f441>0)
                f443 = 0;
        if(f474>0)
                f17 = 0;
        if(f475>0)
                f476 = 0;
        if(f477>0)
                f478 = 0;
        if(f479>0)
                f480 = 0;
        if(f481>0)
                f483 = 0;
        if(f482>0)
                f483 = 0;
        if(f484>0)
                f485 = 0;
        if(f486>0)
                f487 = 0;
        if(f486>0)
                f488 = 0;
        tf = (f0>0)?1:(f1>0)?2:(f2>0)?3:(f3>0)?4:(f4>0)?5:(f5>0)?6:(f6>0)?7:(f7>0)?8:(f8>0)?9:(f9>0)?10:(f10>0)?11:(f11>0)?12:(f12>0)?13:(f13>0)?14:(f14>0)?15:(f15>0)?16:(f16>0)?17:(f17>0)?18:(f18>0)?19:(f19>0)?20:(f20>0)?21:(f21>0)?22:(f22>0)?23:(f23>0)?24:(f24>0)?25:(f25>0)?26:(f26>0)?27:(f27>0)?28:(f28>0)?29:(f29>0)?30:(f30>0)?31:(f31>0)?32:(f32>0)?33:(f33>0)?34:(f34>0)?35:(f35>0)?36:(f36>0)?37:(f37>0)?38:(f38>0)?39:(f39>0)?40:(f40>0)?41:(f41>0)?42:(f42>0)?43:(f43>0)?44:(f44>0)?45:(f45>0)?46:(f46>0)?47:(f47>0)?48:(f48>0)?49:(f49>0)?50:(f50>0)?51:(f51>0)?52:(f52>0)?53:(f53>0)?54:(f54>0)?55:(f55>0)?56:(f56>0)?57:(f57>0)?58:(f58>0)?59:(f59>0)?60:(f60>0)?61:(f61>0)?62:(f62>0)?63:(f63>0)?64:(f64>0)?65:(f65>0)?66:(f66>0)?67:(f67>0)?68:(f68>0)?69:(f69>0)?70:(f70>0)?71:(f71>0)?72:(f72>0)?73:(f73>0)?74:(f74>0)?75:(f75>0)?76:(f76>0)?77:(f77>0)?78:(f78>0)?79:(f79>0)?80:(f80>0)?81:(f81>0)?82:(f82>0)?83:(f83>0)?84:(f84>0)?85:(f85>0)?86:(f86>0)?87:(f87>0)?88:(f88>0)?89:(f89>0)?90:(f90>0)?91:(f91>0)?92:(f92>0)?93:(f93>0)?94:(f94>0)?95:(f95>0)?96:(f96>0)?97:(f97>0)?98:(f98>0)?99:(f99>0)?100:(f100>0)?101:(f101>0)?102:(f102>0)?103:(f103>0)?104:(f104>0)?105:(f105>0)?106:(f106>0)?107:(f107>0)?108:(f108>0)?109:(f109>0)?110:(f110>0)?111:(f111>0)?112:(f112>0)?113:(f113>0)?114:(f114>0)?115:(f115>0)?116:(f116>0)?117:(f117>0)?118:(f118>0)?119:(f119>0)?120:(f120>0)?121:(f121>0)?122:(f122>0)?123:(f123>0)?124:(f124>0)?125:(f125>0)?126:(f126>0)?127:(f127>0)?128:(f128>0)?129:(f129>0)?130:(f130>0)?131:(f131>0)?132:(f132>0)?133:(f133>0)?134:(f134>0)?135:(f135>0)?136:(f136>0)?137:(f137>0)?138:(f138>0)?139:(f139>0)?140:(f140>0)?141:(f141>0)?142:(f142>0)?143:(f143>0)?144:(f144>0)?145:(f145>0)?146:(f146>0)?147:(f147>0)?148:(f148>0)?149:(f149>0)?150:(f150>0)?151:(f151>0)?152:(f152>0)?153:(f153>0)?154:(f154>0)?155:(f155>0)?156:(f156>0)?157:(f157>0)?158:(f158>0)?159:(f159>0)?160:(f160>0)?161:(f161>0)?162:(f162>0)?163:(f163>0)?164:(f164>0)?165:(f165>0)?166:(f166>0)?167:(f167>0)?168:(f168>0)?169:(f169>0)?170:(f170>0)?171:(f171>0)?172:(f172>0)?173:(f173>0)?174:(f174>0)?175:(f175>0)?176:(f176>0)?177:(f177>0)?178:(f178>0)?179:(f179>0)?180:(f180>0)?181:(f181>0)?182:(f182>0)?183:(f183>0)?184:(f184>0)?185:(f185>0)?186:(f186>0)?187:(f187>0)?188:(f188>0)?189:(f189>0)?190:(f190>0)?191:(f191>0)?192:(f192>0)?193:(f193>0)?194:(f194>0)?195:(f195>0)?196:(f196>0)?197:(f197>0)?198:(f198>0)?199:(f199>0)?200:(f200>0)?201:(f201>0)?202:(f202>0)?203:(f203>0)?204:(f204>0)?205:(f205>0)?206:(f206>0)?207:(f207>0)?208:(f208>0)?209:(f209>0)?210:(f210>0)?211:(f211>0)?212:(f212>0)?213:(f213>0)?214:(f214>0)?215:(f215>0)?216:(f216>0)?217:(f217>0)?218:(f218>0)?219:(f219>0)?220:(f220>0)?221:(f221>0)?222:(f222>0)?223:(f223>0)?224:(f224>0)?225:(f225>0)?226:(f226>0)?227:(f227>0)?228:(f228>0)?229:(f229>0)?230:(f230>0)?231:(f231>0)?232:(f232>0)?233:(f233>0)?234:(f234>0)?235:(f235>0)?236:(f236>0)?237:(f237>0)?238:(f238>0)?239:(f239>0)?240:(f240>0)?241:(f241>0)?242:(f242>0)?243:(f243>0)?244:(f244>0)?245:(f245>0)?246:(f246>0)?247:(f247>0)?248:(f248>0)?249:(f249>0)?250:(f250>0)?251:(f251>0)?252:(f252>0)?253:(f253>0)?254:(f254>0)?255:(f255>0)?256:(f256>0)?257:(f257>0)?258:(f258>0)?259:(f259>0)?260:(f260>0)?261:(f261>0)?262:(f262>0)?263:(f263>0)?264:(f264>0)?265:(f265>0)?266:(f266>0)?267:(f267>0)?268:(f268>0)?269:(f269>0)?270:(f270>0)?271:(f271>0)?272:(f272>0)?273:(f273>0)?274:(f274>0)?275:(f275>0)?276:(f276>0)?277:(f277>0)?278:(f278>0)?279:(f279>0)?280:(f280>0)?281:(f281>0)?282:(f282>0)?283:(f283>0)?284:(f284>0)?285:(f285>0)?286:(f286>0)?287:(f287>0)?288:(f288>0)?289:(f289>0)?290:(f290>0)?291:(f291>0)?292:(f292>0)?293:(f293>0)?294:(f294>0)?295:(f295>0)?296:(f296>0)?297:(f297>0)?298:(f298>0)?299:(f299>0)?300:(f300>0)?301:(f301>0)?302:(f302>0)?303:(f303>0)?304:(f304>0)?305:(f305>0)?306:(f306>0)?307:(f307>0)?308:(f308>0)?309:(f309>0)?310:(f310>0)?311:(f311>0)?312:(f312>0)?313:(f313>0)?314:(f314>0)?315:(f315>0)?316:(f316>0)?317:(f317>0)?318:(f318>0)?319:(f319>0)?320:(f320>0)?321:(f321>0)?322:(f322>0)?323:(f323>0)?324:(f324>0)?325:(f325>0)?326:(f326>0)?327:(f327>0)?328:(f328>0)?329:(f329>0)?330:(f330>0)?331:(f331>0)?332:(f332>0)?333:(f333>0)?334:(f334>0)?335:(f335>0)?336:(f336>0)?337:(f337>0)?338:(f338>0)?339:(f339>0)?340:(f340>0)?341:(f341>0)?342:(f342>0)?343:(f343>0)?344:(f344>0)?345:(f345>0)?346:(f346>0)?347:(f347>0)?348:(f348>0)?349:(f349>0)?350:(f350>0)?351:(f351>0)?352:(f352>0)?353:(f353>0)?354:(f354>0)?355:(f355>0)?356:(f356>0)?357:(f357>0)?358:(f358>0)?359:(f359>0)?360:(f360>0)?361:(f361>0)?362:(f362>0)?363:(f363>0)?364:(f364>0)?365:(f365>0)?366:(f366>0)?367:(f367>0)?368:(f368>0)?369:(f369>0)?370:(f370>0)?371:(f371>0)?372:(f372>0)?373:(f373>0)?374:(f374>0)?375:(f375>0)?376:(f376>0)?377:(f377>0)?378:(f378>0)?379:(f379>0)?380:(f380>0)?381:(f381>0)?382:(f382>0)?383:(f383>0)?384:(f384>0)?385:(f385>0)?386:(f386>0)?387:(f387>0)?388:(f388>0)?389:(f389>0)?390:(f390>0)?391:(f391>0)?392:(f392>0)?393:(f393>0)?394:(f394>0)?395:(f395>0)?396:(f396>0)?397:(f397>0)?398:(f398>0)?399:(f399>0)?400:(f400>0)?401:(f401>0)?402:(f402>0)?403:(f403>0)?404:(f404>0)?405:(f405>0)?406:(f406>0)?407:(f407>0)?408:(f408>0)?409:(f409>0)?410:(f410>0)?411:(f411>0)?412:(f412>0)?413:(f413>0)?414:(f414>0)?415:(f415>0)?416:(f416>0)?417:(f417>0)?418:(f418>0)?419:(f419>0)?420:(f420>0)?421:(f421>0)?422:(f422>0)?423:(f423>0)?424:(f424>0)?425:(f425>0)?426:(f426>0)?427:(f427>0)?428:(f428>0)?429:(f429>0)?430:(f430>0)?431:(f431>0)?432:(f432>0)?433:(f433>0)?434:(f434>0)?435:(f435>0)?436:(f436>0)?437:(f437>0)?438:(f438>0)?439:(f439>0)?440:(f440>0)?441:(f441>0)?442:(f442>0)?443:(f443>0)?444:(f444>0)?445:(f445>0)?446:(f446>0)?447:(f447>0)?448:(f448>0)?449:(f449>0)?450:(f450>0)?451:(f451>0)?452:(f452>0)?453:(f453>0)?454:(f454>0)?455:(f455>0)?456:(f456>0)?457:(f457>0)?458:(f458>0)?459:(f459>0)?460:(f460>0)?461:(f461>0)?462:(f462>0)?463:(f463>0)?464:(f464>0)?465:(f465>0)?466:(f466>0)?467:(f467>0)?468:(f468>0)?469:(f469>0)?470:(f470>0)?471:(f471>0)?472:(f472>0)?473:(f473>0)?474:(f474>0)?475:(f475>0)?476:(f476>0)?477:(f477>0)?478:(f478>0)?479:(f479>0)?480:(f480>0)?481:(f481>0)?482:(f482>0)?483:(f483>0)?484:(f484>0)?485:(f485>0)?486:(f486>0)?487:(f487>0)?488:(f488>0)?489:(f489>0)?490:(f490>0)?491:(f491>0)?492:(f492>0)?493:(f493>0)?494:(f494>0)?495:(f495>0)?496:(f496>0)?497:(f497>0)?498:(f498>0)?499:(f499>0)?500:(f500>0)?501:(f501>0)?502:(f502>0)?503:(f503>0)?504:(f504>0)?505:(f505>0)?506:(f506>0)?507:(f507>0)?508:(f508>0)?509:(f509>0)?510:(f510>0)?511:(f511>0)?512:(f512>0)?513:(f513>0)?514:(f514>0)?515:(f515>0)?516:(f516>0)?517:(f517>0)?518:(f518>0)?519:(f519>0)?520:(f520>0)?521:(f521>0)?522:(f522>0)?523:(f523>0)?524:(f524>0)?525:(f525>0)?526:(f526>0)?527:(f527>0)?528:(f528>0)?529:(f529>0)?530:(f530>0)?531:(f531>0)?532:(f532>0)?533:(f533>0)?534:(f534>0)?535:0;
        case(tf)
                1: begin
                        tc = f0;
                        p67 = p67 - tc;
                        p64 = p64 + tc;
                end
                2: begin
                        tc = f1;
                        p91 = p91 - tc;
                        p88 = p88 + tc;
                end
                3: begin
                        tc = f2;
                        p115 = p115 - tc;
                        p112 = p112 + tc;
                end
                4: begin
                        tc = f3;
                        p139 = p139 - tc;
                        p136 = p136 + tc;
                end
                5: begin
                        tc = f4;
                        p163 = p163 - tc;
                        p160 = p160 + tc;
                end
                6: begin
                        tc = f5;
                        p187 = p187 - tc;
                        p184 = p184 + tc;
                end
                7: begin
                        tc = f6;
                        p211 = p211 - tc;
                        p208 = p208 + tc;
                end
                8: begin
                        tc = f7;
                        p235 = p235 - tc;
                        p232 = p232 + tc;
                end
                9: begin
                        tc = f8;
                        p259 = p259 - tc;
                        p256 = p256 + tc;
                end
                10: begin
                        tc = f9;
                        p278 = p278 - tc;
                        p280 = p280 + tc;
                end
                11: begin
                        tc = f10;
                        p297 = p297 - tc;
                        p294 = p294 + tc;
                end
                12: begin
                        tc = f11;
                        p321 = p321 - tc;
                        p318 = p318 + tc;
                end
                13: begin
                        tc = f12;
                        p345 = p345 - tc;
                        p342 = p342 + tc;
                end
                14: begin
                        tc = f13;
                        p364 = p364 - tc;
                        p366 = p366 + tc;
                end
                15: begin
                        tc = f14;
                        p383 = p383 - tc;
                        p380 = p380 + tc;
                end
                16: begin
                        tc = f15;
                        p407 = p407 - tc;
                        p404 = p404 + tc;
                end
                17: begin
                        tc = f16;
                        p426 = p426 - tc;
                        p428 = p428 + tc;
                end
                18: begin
                        tc = f17;
                        p445 = p445 - tc;
                        p442 = p442 + tc;
                end
                19: begin
                        tc = f18;
                        p464 = p464 - tc;
                        p466 = p466 + tc;
                end
                20: begin
                        tc = f19;
                        p478 = p478 - tc;
                        p480 = p480 + tc;
                end
                21: begin
                        tc = f20;
                        p68 = p68 - tc;
                        p64 = p64 + tc;
                end
                22: begin
                        tc = f21;
                        p62 = p62 - tc;
                end
                23: begin
                        tc = f22;
                        p66 = p66 - tc;
                        p68 = p68 + tc;
                end
                24: begin
                        tc = f23;
                        p63 = p63 - tc*2;
                        p69 = p69 + tc;
                end
                25: begin
                        tc = f24;
                        p70 = p70 - tc;
                        p67 = p67 + tc;
                end
                26: begin
                        tc = f25;
                        p63 = p63 - tc;
                        p72 = p72 - tc;
                        p71 = p71 + tc;
                end
                27: begin
                        tc = f26;
                        p73 = p73 - tc;
                        p70 = p70 + tc;
                end
                28: begin
                        tc = f27;
                        p62 = p62 - tc;
                        p65 = p65 + tc;
                        p74 = p74 + tc;
                end
                29: begin
                        tc = f28;
                        p62 = p62 - tc;
                        p74 = p74 + tc;
                end
                30: begin
                        tc = f29;
                        p75 = p75 - tc;
                        p73 = p73 + tc;
                end
                31: begin
                        tc = f30;
                        p69 = p69 - tc;
                        p63 = p63 + tc;
                end
                32: begin
                        tc = f31;
                        p76 = p76 - tc;
                        p75 = p75 + tc;
                end
                33: begin
                        tc = f32;
                        p74 = p74 - tc;
                        p62 = p62 + tc*2;
                end
                34: begin
                        tc = f33;
                        p64 = p64 - tc;
                        p71 = p71 - tc;
                        p72 = p72 + tc;
                        p76 = p76 + tc;
                end
                35: begin
                        tc = f34;
                        p64 = p64 - tc;
                        p76 = p76 + tc;
                end
                36: begin
                        tc = f35;
                        p21 = p21 - tc;
                        p62 = p62 + tc;
                        p77 = p77 + tc;
                end
                37: begin
                        tc = f36;
                        p77 = p77 - tc;
                        p21 = p21 + tc;
                end
                38: begin
                        tc = f37;
                        p79 = p79 - tc;
                        p78 = p78 + tc;
                end
                39: begin
                        tc = f38;
                        p80 = p80 - tc;
                        p79 = p79 + tc;
                end
                40: begin
                        tc = f39;
                        p22 = p22 - tc;
                        p63 = p63 + tc;
                        p81 = p81 + tc;
                end
                41: begin
                        tc = f40;
                        p81 = p81 - tc;
                        p22 = p22 + tc;
                end
                42: begin
                        tc = f41;
                        p83 = p83 - tc;
                        p82 = p82 + tc;
                end
                43: begin
                        tc = f42;
                        p84 = p84 - tc;
                        p83 = p83 + tc;
                end
                44: begin
                        tc = f43;
                        p78 = p78 - tc;
                        p82 = p82 - tc;
                        p0 = p0 + tc;
                end
                45: begin
                        tc = f44;
                        p64 = p64 - tc;
                        p80 = p80 + tc;
                        p84 = p84 + tc;
                end
                46: begin
                        tc = f45;
                        p65 = p65 - tc;
                        p23 = p23 + tc;
                end
                47: begin
                        tc = f46;
                        p23 = p23 - tc;
                end
                48: begin
                        tc = f47;
                        p85 = p85 - tc;
                        p66 = p66 + tc;
                end
                49: begin
                        tc = f48;
                        p1 = p1 - tc;
                        p85 = p85 + tc;
                end
                50: begin
                        tc = f49;
                        p92 = p92 - tc;
                        p88 = p88 + tc;
                end
                51: begin
                        tc = f50;
                        p86 = p86 - tc;
                end
                52: begin
                        tc = f51;
                        p90 = p90 - tc;
                        p92 = p92 + tc;
                end
                53: begin
                        tc = f52;
                        p87 = p87 - tc*2;
                        p93 = p93 + tc;
                end
                54: begin
                        tc = f53;
                        p94 = p94 - tc;
                        p91 = p91 + tc;
                end
                55: begin
                        tc = f54;
                        p87 = p87 - tc;
                        p96 = p96 - tc;
                        p95 = p95 + tc;
                end
                56: begin
                        tc = f55;
                        p97 = p97 - tc;
                        p94 = p94 + tc;
                end
                57: begin
                        tc = f56;
                        p86 = p86 - tc;
                        p89 = p89 + tc;
                        p98 = p98 + tc;
                end
                58: begin
                        tc = f57;
                        p86 = p86 - tc;
                        p98 = p98 + tc;
                end
                59: begin
                        tc = f58;
                        p99 = p99 - tc;
                        p97 = p97 + tc;
                end
                60: begin
                        tc = f59;
                        p93 = p93 - tc;
                        p87 = p87 + tc;
                end
                61: begin
                        tc = f60;
                        p100 = p100 - tc;
                        p99 = p99 + tc;
                end
                62: begin
                        tc = f61;
                        p98 = p98 - tc;
                        p86 = p86 + tc*2;
                end
                63: begin
                        tc = f62;
                        p88 = p88 - tc;
                        p95 = p95 - tc;
                        p96 = p96 + tc;
                        p100 = p100 + tc;
                end
                64: begin
                        tc = f63;
                        p88 = p88 - tc;
                        p100 = p100 + tc;
                end
                65: begin
                        tc = f64;
                        p23 = p23 - tc;
                        p86 = p86 + tc;
                        p101 = p101 + tc;
                end
                66: begin
                        tc = f65;
                        p101 = p101 - tc;
                        p23 = p23 + tc;
                end
                67: begin
                        tc = f66;
                        p103 = p103 - tc;
                        p102 = p102 + tc;
                end
                68: begin
                        tc = f67;
                        p104 = p104 - tc;
                        p103 = p103 + tc;
                end
                69: begin
                        tc = f68;
                        p24 = p24 - tc;
                        p87 = p87 + tc;
                        p105 = p105 + tc;
                end
                70: begin
                        tc = f69;
                        p105 = p105 - tc;
                        p24 = p24 + tc;
                end
                71: begin
                        tc = f70;
                        p107 = p107 - tc;
                        p106 = p106 + tc;
                end
                72: begin
                        tc = f71;
                        p108 = p108 - tc;
                        p107 = p107 + tc;
                end
                73: begin
                        tc = f72;
                        p102 = p102 - tc;
                        p106 = p106 - tc;
                        p1 = p1 + tc;
                end
                74: begin
                        tc = f73;
                        p88 = p88 - tc;
                        p104 = p104 + tc;
                        p108 = p108 + tc;
                end
                75: begin
                        tc = f74;
                        p89 = p89 - tc;
                        p25 = p25 + tc;
                end
                76: begin
                        tc = f75;
                        p25 = p25 - tc;
                end
                77: begin
                        tc = f76;
                        p109 = p109 - tc;
                        p90 = p90 + tc;
                end
                78: begin
                        tc = f77;
                        p2 = p2 - tc;
                        p109 = p109 + tc;
                end
                79: begin
                        tc = f78;
                        p116 = p116 - tc;
                        p112 = p112 + tc;
                end
                80: begin
                        tc = f79;
                        p110 = p110 - tc;
                end
                81: begin
                        tc = f80;
                        p114 = p114 - tc;
                        p116 = p116 + tc;
                end
                82: begin
                        tc = f81;
                        p111 = p111 - tc*2;
                        p117 = p117 + tc;
                end
                83: begin
                        tc = f82;
                        p118 = p118 - tc;
                        p115 = p115 + tc;
                end
                84: begin
                        tc = f83;
                        p111 = p111 - tc;
                        p120 = p120 - tc;
                        p119 = p119 + tc;
                end
                85: begin
                        tc = f84;
                        p121 = p121 - tc;
                        p118 = p118 + tc;
                end
                86: begin
                        tc = f85;
                        p110 = p110 - tc;
                        p113 = p113 + tc;
                        p122 = p122 + tc;
                end
                87: begin
                        tc = f86;
                        p110 = p110 - tc;
                        p122 = p122 + tc;
                end
                88: begin
                        tc = f87;
                        p123 = p123 - tc;
                        p121 = p121 + tc;
                end
                89: begin
                        tc = f88;
                        p117 = p117 - tc;
                        p111 = p111 + tc;
                end
                90: begin
                        tc = f89;
                        p124 = p124 - tc;
                        p123 = p123 + tc;
                end
                91: begin
                        tc = f90;
                        p122 = p122 - tc;
                        p110 = p110 + tc*2;
                end
                92: begin
                        tc = f91;
                        p112 = p112 - tc;
                        p119 = p119 - tc;
                        p120 = p120 + tc;
                        p124 = p124 + tc;
                end
                93: begin
                        tc = f92;
                        p112 = p112 - tc;
                        p124 = p124 + tc;
                end
                94: begin
                        tc = f93;
                        p25 = p25 - tc;
                        p110 = p110 + tc;
                        p125 = p125 + tc;
                end
                95: begin
                        tc = f94;
                        p125 = p125 - tc;
                        p25 = p25 + tc;
                end
                96: begin
                        tc = f95;
                        p127 = p127 - tc;
                        p126 = p126 + tc;
                end
                97: begin
                        tc = f96;
                        p128 = p128 - tc;
                        p127 = p127 + tc;
                end
                98: begin
                        tc = f97;
                        p26 = p26 - tc;
                        p111 = p111 + tc;
                        p129 = p129 + tc;
                end
                99: begin
                        tc = f98;
                        p129 = p129 - tc;
                        p26 = p26 + tc;
                end
                100: begin
                        tc = f99;
                        p131 = p131 - tc;
                        p130 = p130 + tc;
                end
                101: begin
                        tc = f100;
                        p132 = p132 - tc;
                        p131 = p131 + tc;
                end
                102: begin
                        tc = f101;
                        p126 = p126 - tc;
                        p130 = p130 - tc;
                        p2 = p2 + tc;
                end
                103: begin
                        tc = f102;
                        p112 = p112 - tc;
                        p128 = p128 + tc;
                        p132 = p132 + tc;
                end
                104: begin
                        tc = f103;
                        p113 = p113 - tc;
                        p27 = p27 + tc;
                end
                105: begin
                        tc = f104;
                        p27 = p27 - tc;
                end
                106: begin
                        tc = f105;
                        p133 = p133 - tc;
                        p114 = p114 + tc;
                end
                107: begin
                        tc = f106;
                        p3 = p3 - tc;
                        p133 = p133 + tc;
                end
                108: begin
                        tc = f107;
                        p140 = p140 - tc;
                        p136 = p136 + tc;
                end
                109: begin
                        tc = f108;
                        p134 = p134 - tc;
                end
                110: begin
                        tc = f109;
                        p138 = p138 - tc;
                        p140 = p140 + tc;
                end
                111: begin
                        tc = f110;
                        p135 = p135 - tc*2;
                        p141 = p141 + tc;
                end
                112: begin
                        tc = f111;
                        p142 = p142 - tc;
                        p139 = p139 + tc;
                end
                113: begin
                        tc = f112;
                        p135 = p135 - tc;
                        p144 = p144 - tc;
                        p143 = p143 + tc;
                end
                114: begin
                        tc = f113;
                        p145 = p145 - tc;
                        p142 = p142 + tc;
                end
                115: begin
                        tc = f114;
                        p134 = p134 - tc;
                        p137 = p137 + tc;
                        p146 = p146 + tc;
                end
                116: begin
                        tc = f115;
                        p134 = p134 - tc;
                        p146 = p146 + tc;
                end
                117: begin
                        tc = f116;
                        p147 = p147 - tc;
                        p145 = p145 + tc;
                end
                118: begin
                        tc = f117;
                        p141 = p141 - tc;
                        p135 = p135 + tc;
                end
                119: begin
                        tc = f118;
                        p148 = p148 - tc;
                        p147 = p147 + tc;
                end
                120: begin
                        tc = f119;
                        p146 = p146 - tc;
                        p134 = p134 + tc*2;
                end
                121: begin
                        tc = f120;
                        p136 = p136 - tc;
                        p143 = p143 - tc;
                        p144 = p144 + tc;
                        p148 = p148 + tc;
                end
                122: begin
                        tc = f121;
                        p136 = p136 - tc;
                        p148 = p148 + tc;
                end
                123: begin
                        tc = f122;
                        p27 = p27 - tc;
                        p134 = p134 + tc;
                        p149 = p149 + tc;
                end
                124: begin
                        tc = f123;
                        p149 = p149 - tc;
                        p27 = p27 + tc;
                end
                125: begin
                        tc = f124;
                        p151 = p151 - tc;
                        p150 = p150 + tc;
                end
                126: begin
                        tc = f125;
                        p152 = p152 - tc;
                        p151 = p151 + tc;
                end
                127: begin
                        tc = f126;
                        p28 = p28 - tc;
                        p135 = p135 + tc;
                        p153 = p153 + tc;
                end
                128: begin
                        tc = f127;
                        p153 = p153 - tc;
                        p28 = p28 + tc;
                end
                129: begin
                        tc = f128;
                        p155 = p155 - tc;
                        p154 = p154 + tc;
                end
                130: begin
                        tc = f129;
                        p156 = p156 - tc;
                        p155 = p155 + tc;
                end
                131: begin
                        tc = f130;
                        p150 = p150 - tc;
                        p154 = p154 - tc;
                        p3 = p3 + tc;
                end
                132: begin
                        tc = f131;
                        p136 = p136 - tc;
                        p152 = p152 + tc;
                        p156 = p156 + tc;
                end
                133: begin
                        tc = f132;
                        p137 = p137 - tc;
                        p29 = p29 + tc;
                end
                134: begin
                        tc = f133;
                        p29 = p29 - tc;
                end
                135: begin
                        tc = f134;
                        p157 = p157 - tc;
                        p138 = p138 + tc;
                end
                136: begin
                        tc = f135;
                        p4 = p4 - tc;
                        p157 = p157 + tc;
                end
                137: begin
                        tc = f136;
                        p164 = p164 - tc;
                        p160 = p160 + tc;
                end
                138: begin
                        tc = f137;
                        p158 = p158 - tc;
                end
                139: begin
                        tc = f138;
                        p162 = p162 - tc;
                        p164 = p164 + tc;
                end
                140: begin
                        tc = f139;
                        p159 = p159 - tc*2;
                        p165 = p165 + tc;
                end
                141: begin
                        tc = f140;
                        p166 = p166 - tc;
                        p163 = p163 + tc;
                end
                142: begin
                        tc = f141;
                        p159 = p159 - tc;
                        p168 = p168 - tc;
                        p167 = p167 + tc;
                end
                143: begin
                        tc = f142;
                        p169 = p169 - tc;
                        p166 = p166 + tc;
                end
                144: begin
                        tc = f143;
                        p158 = p158 - tc;
                        p161 = p161 + tc;
                        p170 = p170 + tc;
                end
                145: begin
                        tc = f144;
                        p158 = p158 - tc;
                        p170 = p170 + tc;
                end
                146: begin
                        tc = f145;
                        p171 = p171 - tc;
                        p169 = p169 + tc;
                end
                147: begin
                        tc = f146;
                        p165 = p165 - tc;
                        p159 = p159 + tc;
                end
                148: begin
                        tc = f147;
                        p172 = p172 - tc;
                        p171 = p171 + tc;
                end
                149: begin
                        tc = f148;
                        p170 = p170 - tc;
                        p158 = p158 + tc*2;
                end
                150: begin
                        tc = f149;
                        p160 = p160 - tc;
                        p167 = p167 - tc;
                        p168 = p168 + tc;
                        p172 = p172 + tc;
                end
                151: begin
                        tc = f150;
                        p160 = p160 - tc;
                        p172 = p172 + tc;
                end
                152: begin
                        tc = f151;
                        p29 = p29 - tc;
                        p158 = p158 + tc;
                        p173 = p173 + tc;
                end
                153: begin
                        tc = f152;
                        p173 = p173 - tc;
                        p29 = p29 + tc;
                end
                154: begin
                        tc = f153;
                        p175 = p175 - tc;
                        p174 = p174 + tc;
                end
                155: begin
                        tc = f154;
                        p176 = p176 - tc;
                        p175 = p175 + tc;
                end
                156: begin
                        tc = f155;
                        p30 = p30 - tc;
                        p159 = p159 + tc;
                        p177 = p177 + tc;
                end
                157: begin
                        tc = f156;
                        p177 = p177 - tc;
                        p30 = p30 + tc;
                end
                158: begin
                        tc = f157;
                        p179 = p179 - tc;
                        p178 = p178 + tc;
                end
                159: begin
                        tc = f158;
                        p180 = p180 - tc;
                        p179 = p179 + tc;
                end
                160: begin
                        tc = f159;
                        p174 = p174 - tc;
                        p178 = p178 - tc;
                        p4 = p4 + tc;
                end
                161: begin
                        tc = f160;
                        p160 = p160 - tc;
                        p176 = p176 + tc;
                        p180 = p180 + tc;
                end
                162: begin
                        tc = f161;
                        p161 = p161 - tc;
                        p31 = p31 + tc;
                end
                163: begin
                        tc = f162;
                        p31 = p31 - tc;
                end
                164: begin
                        tc = f163;
                        p181 = p181 - tc;
                        p162 = p162 + tc;
                end
                165: begin
                        tc = f164;
                        p5 = p5 - tc;
                        p181 = p181 + tc;
                end
                166: begin
                        tc = f165;
                        p188 = p188 - tc;
                        p184 = p184 + tc;
                end
                167: begin
                        tc = f166;
                        p182 = p182 - tc;
                end
                168: begin
                        tc = f167;
                        p186 = p186 - tc;
                        p188 = p188 + tc;
                end
                169: begin
                        tc = f168;
                        p183 = p183 - tc*2;
                        p189 = p189 + tc;
                end
                170: begin
                        tc = f169;
                        p190 = p190 - tc;
                        p187 = p187 + tc;
                end
                171: begin
                        tc = f170;
                        p183 = p183 - tc;
                        p192 = p192 - tc;
                        p191 = p191 + tc;
                end
                172: begin
                        tc = f171;
                        p193 = p193 - tc;
                        p190 = p190 + tc;
                end
                173: begin
                        tc = f172;
                        p182 = p182 - tc;
                        p185 = p185 + tc;
                        p194 = p194 + tc;
                end
                174: begin
                        tc = f173;
                        p182 = p182 - tc;
                        p194 = p194 + tc;
                end
                175: begin
                        tc = f174;
                        p195 = p195 - tc;
                        p193 = p193 + tc;
                end
                176: begin
                        tc = f175;
                        p189 = p189 - tc;
                        p183 = p183 + tc;
                end
                177: begin
                        tc = f176;
                        p196 = p196 - tc;
                        p195 = p195 + tc;
                end
                178: begin
                        tc = f177;
                        p194 = p194 - tc;
                        p182 = p182 + tc*2;
                end
                179: begin
                        tc = f178;
                        p184 = p184 - tc;
                        p191 = p191 - tc;
                        p192 = p192 + tc;
                        p196 = p196 + tc;
                end
                180: begin
                        tc = f179;
                        p184 = p184 - tc;
                        p196 = p196 + tc;
                end
                181: begin
                        tc = f180;
                        p32 = p32 - tc;
                        p182 = p182 + tc;
                        p197 = p197 + tc;
                end
                182: begin
                        tc = f181;
                        p197 = p197 - tc;
                        p32 = p32 + tc;
                end
                183: begin
                        tc = f182;
                        p199 = p199 - tc;
                        p198 = p198 + tc;
                end
                184: begin
                        tc = f183;
                        p200 = p200 - tc;
                        p199 = p199 + tc;
                end
                185: begin
                        tc = f184;
                        p33 = p33 - tc;
                        p183 = p183 + tc;
                        p201 = p201 + tc;
                end
                186: begin
                        tc = f185;
                        p201 = p201 - tc;
                        p33 = p33 + tc;
                end
                187: begin
                        tc = f186;
                        p203 = p203 - tc;
                        p202 = p202 + tc;
                end
                188: begin
                        tc = f187;
                        p204 = p204 - tc;
                        p203 = p203 + tc;
                end
                189: begin
                        tc = f188;
                        p198 = p198 - tc;
                        p202 = p202 - tc;
                        p5 = p5 + tc;
                end
                190: begin
                        tc = f189;
                        p184 = p184 - tc;
                        p200 = p200 + tc;
                        p204 = p204 + tc;
                end
                191: begin
                        tc = f190;
                        p185 = p185 - tc;
                        p34 = p34 + tc;
                end
                192: begin
                        tc = f191;
                        p34 = p34 - tc;
                end
                193: begin
                        tc = f192;
                        p205 = p205 - tc;
                        p186 = p186 + tc;
                end
                194: begin
                        tc = f193;
                        p6 = p6 - tc;
                        p205 = p205 + tc;
                end
                195: begin
                        tc = f194;
                        p212 = p212 - tc;
                        p208 = p208 + tc;
                end
                196: begin
                        tc = f195;
                        p206 = p206 - tc;
                end
                197: begin
                        tc = f196;
                        p210 = p210 - tc;
                        p212 = p212 + tc;
                end
                198: begin
                        tc = f197;
                        p207 = p207 - tc*2;
                        p213 = p213 + tc;
                end
                199: begin
                        tc = f198;
                        p214 = p214 - tc;
                        p211 = p211 + tc;
                end
                200: begin
                        tc = f199;
                        p207 = p207 - tc;
                        p216 = p216 - tc;
                        p215 = p215 + tc;
                end
                201: begin
                        tc = f200;
                        p217 = p217 - tc;
                        p214 = p214 + tc;
                end
                202: begin
                        tc = f201;
                        p206 = p206 - tc;
                        p209 = p209 + tc;
                        p218 = p218 + tc;
                end
                203: begin
                        tc = f202;
                        p206 = p206 - tc;
                        p218 = p218 + tc;
                end
                204: begin
                        tc = f203;
                        p219 = p219 - tc;
                        p217 = p217 + tc;
                end
                205: begin
                        tc = f204;
                        p213 = p213 - tc;
                        p207 = p207 + tc;
                end
                206: begin
                        tc = f205;
                        p220 = p220 - tc;
                        p219 = p219 + tc;
                end
                207: begin
                        tc = f206;
                        p218 = p218 - tc;
                        p206 = p206 + tc*2;
                end
                208: begin
                        tc = f207;
                        p208 = p208 - tc;
                        p215 = p215 - tc;
                        p216 = p216 + tc;
                        p220 = p220 + tc;
                end
                209: begin
                        tc = f208;
                        p208 = p208 - tc;
                        p220 = p220 + tc;
                end
                210: begin
                        tc = f209;
                        p34 = p34 - tc;
                        p206 = p206 + tc;
                        p221 = p221 + tc;
                end
                211: begin
                        tc = f210;
                        p221 = p221 - tc;
                        p34 = p34 + tc;
                end
                212: begin
                        tc = f211;
                        p223 = p223 - tc;
                        p222 = p222 + tc;
                end
                213: begin
                        tc = f212;
                        p224 = p224 - tc;
                        p223 = p223 + tc;
                end
                214: begin
                        tc = f213;
                        p35 = p35 - tc;
                        p207 = p207 + tc;
                        p225 = p225 + tc;
                end
                215: begin
                        tc = f214;
                        p225 = p225 - tc;
                        p35 = p35 + tc;
                end
                216: begin
                        tc = f215;
                        p227 = p227 - tc;
                        p226 = p226 + tc;
                end
                217: begin
                        tc = f216;
                        p228 = p228 - tc;
                        p227 = p227 + tc;
                end
                218: begin
                        tc = f217;
                        p222 = p222 - tc;
                        p226 = p226 - tc;
                        p6 = p6 + tc;
                end
                219: begin
                        tc = f218;
                        p208 = p208 - tc;
                        p224 = p224 + tc;
                        p228 = p228 + tc;
                end
                220: begin
                        tc = f219;
                        p209 = p209 - tc;
                        p36 = p36 + tc;
                end
                221: begin
                        tc = f220;
                        p36 = p36 - tc;
                end
                222: begin
                        tc = f221;
                        p229 = p229 - tc;
                        p210 = p210 + tc;
                end
                223: begin
                        tc = f222;
                        p7 = p7 - tc;
                        p229 = p229 + tc;
                end
                224: begin
                        tc = f223;
                        p236 = p236 - tc;
                        p232 = p232 + tc;
                end
                225: begin
                        tc = f224;
                        p230 = p230 - tc;
                end
                226: begin
                        tc = f225;
                        p234 = p234 - tc;
                        p236 = p236 + tc;
                end
                227: begin
                        tc = f226;
                        p231 = p231 - tc*2;
                        p237 = p237 + tc;
                end
                228: begin
                        tc = f227;
                        p238 = p238 - tc;
                        p235 = p235 + tc;
                end
                229: begin
                        tc = f228;
                        p231 = p231 - tc;
                        p240 = p240 - tc;
                        p239 = p239 + tc;
                end
                230: begin
                        tc = f229;
                        p241 = p241 - tc;
                        p238 = p238 + tc;
                end
                231: begin
                        tc = f230;
                        p230 = p230 - tc;
                        p233 = p233 + tc;
                        p242 = p242 + tc;
                end
                232: begin
                        tc = f231;
                        p230 = p230 - tc;
                        p242 = p242 + tc;
                end
                233: begin
                        tc = f232;
                        p243 = p243 - tc;
                        p241 = p241 + tc;
                end
                234: begin
                        tc = f233;
                        p237 = p237 - tc;
                        p231 = p231 + tc;
                end
                235: begin
                        tc = f234;
                        p244 = p244 - tc;
                        p243 = p243 + tc;
                end
                236: begin
                        tc = f235;
                        p242 = p242 - tc;
                        p230 = p230 + tc*2;
                end
                237: begin
                        tc = f236;
                        p232 = p232 - tc;
                        p239 = p239 - tc;
                        p240 = p240 + tc;
                        p244 = p244 + tc;
                end
                238: begin
                        tc = f237;
                        p232 = p232 - tc;
                        p244 = p244 + tc;
                end
                239: begin
                        tc = f238;
                        p36 = p36 - tc;
                        p230 = p230 + tc;
                        p245 = p245 + tc;
                end
                240: begin
                        tc = f239;
                        p245 = p245 - tc;
                        p36 = p36 + tc;
                end
                241: begin
                        tc = f240;
                        p247 = p247 - tc;
                        p246 = p246 + tc;
                end
                242: begin
                        tc = f241;
                        p248 = p248 - tc;
                        p247 = p247 + tc;
                end
                243: begin
                        tc = f242;
                        p37 = p37 - tc;
                        p231 = p231 + tc;
                        p249 = p249 + tc;
                end
                244: begin
                        tc = f243;
                        p249 = p249 - tc;
                        p37 = p37 + tc;
                end
                245: begin
                        tc = f244;
                        p251 = p251 - tc;
                        p250 = p250 + tc;
                end
                246: begin
                        tc = f245;
                        p252 = p252 - tc;
                        p251 = p251 + tc;
                end
                247: begin
                        tc = f246;
                        p246 = p246 - tc;
                        p250 = p250 - tc;
                        p7 = p7 + tc;
                end
                248: begin
                        tc = f247;
                        p232 = p232 - tc;
                        p248 = p248 + tc;
                        p252 = p252 + tc;
                end
                249: begin
                        tc = f248;
                        p233 = p233 - tc;
                        p38 = p38 + tc;
                end
                250: begin
                        tc = f249;
                        p38 = p38 - tc;
                end
                251: begin
                        tc = f250;
                        p253 = p253 - tc;
                        p234 = p234 + tc;
                end
                252: begin
                        tc = f251;
                        p8 = p8 - tc;
                        p253 = p253 + tc;
                end
                253: begin
                        tc = f252;
                        p260 = p260 - tc;
                        p256 = p256 + tc;
                end
                254: begin
                        tc = f253;
                        p254 = p254 - tc;
                end
                255: begin
                        tc = f254;
                        p258 = p258 - tc;
                        p260 = p260 + tc;
                end
                256: begin
                        tc = f255;
                        p255 = p255 - tc*2;
                        p261 = p261 + tc;
                end
                257: begin
                        tc = f256;
                        p262 = p262 - tc;
                        p259 = p259 + tc;
                end
                258: begin
                        tc = f257;
                        p255 = p255 - tc;
                        p264 = p264 - tc;
                        p263 = p263 + tc;
                end
                259: begin
                        tc = f258;
                        p265 = p265 - tc;
                        p262 = p262 + tc;
                end
                260: begin
                        tc = f259;
                        p254 = p254 - tc;
                        p257 = p257 + tc;
                        p266 = p266 + tc;
                end
                261: begin
                        tc = f260;
                        p254 = p254 - tc;
                        p266 = p266 + tc;
                end
                262: begin
                        tc = f261;
                        p267 = p267 - tc;
                        p265 = p265 + tc;
                end
                263: begin
                        tc = f262;
                        p261 = p261 - tc;
                        p255 = p255 + tc;
                end
                264: begin
                        tc = f263;
                        p268 = p268 - tc;
                        p267 = p267 + tc;
                end
                265: begin
                        tc = f264;
                        p266 = p266 - tc;
                        p254 = p254 + tc*2;
                end
                266: begin
                        tc = f265;
                        p256 = p256 - tc;
                        p263 = p263 - tc;
                        p264 = p264 + tc;
                        p268 = p268 + tc;
                end
                267: begin
                        tc = f266;
                        p256 = p256 - tc;
                        p268 = p268 + tc;
                end
                268: begin
                        tc = f267;
                        p38 = p38 - tc;
                        p254 = p254 + tc;
                        p269 = p269 + tc;
                end
                269: begin
                        tc = f268;
                        p269 = p269 - tc;
                        p38 = p38 + tc;
                end
                270: begin
                        tc = f269;
                        p271 = p271 - tc;
                        p270 = p270 + tc;
                end
                271: begin
                        tc = f270;
                        p272 = p272 - tc;
                        p271 = p271 + tc;
                end
                272: begin
                        tc = f271;
                        p39 = p39 - tc;
                        p255 = p255 + tc;
                        p273 = p273 + tc;
                end
                273: begin
                        tc = f272;
                        p273 = p273 - tc;
                        p39 = p39 + tc;
                end
                274: begin
                        tc = f273;
                        p275 = p275 - tc;
                        p274 = p274 + tc;
                end
                275: begin
                        tc = f274;
                        p276 = p276 - tc;
                        p275 = p275 + tc;
                end
                276: begin
                        tc = f275;
                        p270 = p270 - tc;
                        p274 = p274 - tc;
                        p8 = p8 + tc;
                end
                277: begin
                        tc = f276;
                        p256 = p256 - tc;
                        p272 = p272 + tc;
                        p276 = p276 + tc;
                end
                278: begin
                        tc = f277;
                        p257 = p257 - tc;
                        p40 = p40 + tc;
                end
                279: begin
                        tc = f278;
                        p40 = p40 - tc;
                end
                280: begin
                        tc = f279;
                        p277 = p277 - tc;
                        p258 = p258 + tc;
                end
                281: begin
                        tc = f280;
                        p9 = p9 - tc;
                        p277 = p277 + tc;
                end
                282: begin
                        tc = f281;
                        p279 = p279 - tc;
                        p280 = p280 + tc;
                end
                283: begin
                        tc = f282;
                        p282 = p282 - tc;
                        p281 = p281 + tc;
                end
                284: begin
                        tc = f283;
                        p31 = p31 - tc;
                        p278 = p278 + tc;
                        p283 = p283 + tc;
                end
                285: begin
                        tc = f284;
                        p283 = p283 - tc;
                        p31 = p31 + tc;
                end
                286: begin
                        tc = f285;
                        p285 = p285 - tc;
                        p284 = p284 + tc;
                end
                287: begin
                        tc = f286;
                        p286 = p286 - tc;
                        p285 = p285 + tc;
                end
                288: begin
                        tc = f287;
                        p40 = p40 - tc;
                        p279 = p279 + tc;
                        p287 = p287 + tc;
                end
                289: begin
                        tc = f288;
                        p287 = p287 - tc;
                        p40 = p40 + tc;
                end
                290: begin
                        tc = f289;
                        p289 = p289 - tc;
                        p288 = p288 + tc;
                end
                291: begin
                        tc = f290;
                        p290 = p290 - tc;
                        p289 = p289 + tc;
                end
                292: begin
                        tc = f291;
                        p284 = p284 - tc;
                        p288 = p288 - tc;
                        p9 = p9 + tc;
                end
                293: begin
                        tc = f292;
                        p281 = p281 - tc;
                        p286 = p286 + tc;
                        p290 = p290 + tc;
                end
                294: begin
                        tc = f293;
                        p280 = p280 - tc;
                        p41 = p41 + tc;
                end
                295: begin
                        tc = f294;
                        p41 = p41 - tc;
                end
                296: begin
                        tc = f295;
                        p291 = p291 - tc;
                        p282 = p282 + tc;
                end
                297: begin
                        tc = f296;
                        p10 = p10 - tc;
                        p291 = p291 + tc;
                end
                298: begin
                        tc = f297;
                        p298 = p298 - tc;
                        p294 = p294 + tc;
                end
                299: begin
                        tc = f298;
                        p292 = p292 - tc;
                end
                300: begin
                        tc = f299;
                        p296 = p296 - tc;
                        p298 = p298 + tc;
                end
                301: begin
                        tc = f300;
                        p293 = p293 - tc*2;
                        p299 = p299 + tc;
                end
                302: begin
                        tc = f301;
                        p300 = p300 - tc;
                        p297 = p297 + tc;
                end
                303: begin
                        tc = f302;
                        p293 = p293 - tc;
                        p302 = p302 - tc;
                        p301 = p301 + tc;
                end
                304: begin
                        tc = f303;
                        p303 = p303 - tc;
                        p300 = p300 + tc;
                end
                305: begin
                        tc = f304;
                        p292 = p292 - tc;
                        p295 = p295 + tc;
                        p304 = p304 + tc;
                end
                306: begin
                        tc = f305;
                        p292 = p292 - tc;
                        p304 = p304 + tc;
                end
                307: begin
                        tc = f306;
                        p305 = p305 - tc;
                        p303 = p303 + tc;
                end
                308: begin
                        tc = f307;
                        p299 = p299 - tc;
                        p293 = p293 + tc;
                end
                309: begin
                        tc = f308;
                        p306 = p306 - tc;
                        p305 = p305 + tc;
                end
                310: begin
                        tc = f309;
                        p304 = p304 - tc;
                        p292 = p292 + tc*2;
                end
                311: begin
                        tc = f310;
                        p294 = p294 - tc;
                        p301 = p301 - tc;
                        p302 = p302 + tc;
                        p306 = p306 + tc;
                end
                312: begin
                        tc = f311;
                        p294 = p294 - tc;
                        p306 = p306 + tc;
                end
                313: begin
                        tc = f312;
                        p42 = p42 - tc;
                        p292 = p292 + tc;
                        p307 = p307 + tc;
                end
                314: begin
                        tc = f313;
                        p307 = p307 - tc;
                        p42 = p42 + tc;
                end
                315: begin
                        tc = f314;
                        p309 = p309 - tc;
                        p308 = p308 + tc;
                end
                316: begin
                        tc = f315;
                        p310 = p310 - tc;
                        p309 = p309 + tc;
                end
                317: begin
                        tc = f316;
                        p43 = p43 - tc;
                        p293 = p293 + tc;
                        p311 = p311 + tc;
                end
                318: begin
                        tc = f317;
                        p311 = p311 - tc;
                        p43 = p43 + tc;
                end
                319: begin
                        tc = f318;
                        p313 = p313 - tc;
                        p312 = p312 + tc;
                end
                320: begin
                        tc = f319;
                        p314 = p314 - tc;
                        p313 = p313 + tc;
                end
                321: begin
                        tc = f320;
                        p308 = p308 - tc;
                        p312 = p312 - tc;
                        p10 = p10 + tc;
                end
                322: begin
                        tc = f321;
                        p294 = p294 - tc;
                        p310 = p310 + tc;
                        p314 = p314 + tc;
                end
                323: begin
                        tc = f322;
                        p295 = p295 - tc;
                        p44 = p44 + tc;
                end
                324: begin
                        tc = f323;
                        p44 = p44 - tc;
                end
                325: begin
                        tc = f324;
                        p315 = p315 - tc;
                        p296 = p296 + tc;
                end
                326: begin
                        tc = f325;
                        p11 = p11 - tc;
                        p315 = p315 + tc;
                end
                327: begin
                        tc = f326;
                        p322 = p322 - tc;
                        p318 = p318 + tc;
                end
                328: begin
                        tc = f327;
                        p316 = p316 - tc;
                end
                329: begin
                        tc = f328;
                        p320 = p320 - tc;
                        p322 = p322 + tc;
                end
                330: begin
                        tc = f329;
                        p317 = p317 - tc*2;
                        p323 = p323 + tc;
                end
                331: begin
                        tc = f330;
                        p324 = p324 - tc;
                        p321 = p321 + tc;
                end
                332: begin
                        tc = f331;
                        p317 = p317 - tc;
                        p326 = p326 - tc;
                        p325 = p325 + tc;
                end
                333: begin
                        tc = f332;
                        p327 = p327 - tc;
                        p324 = p324 + tc;
                end
                334: begin
                        tc = f333;
                        p316 = p316 - tc;
                        p319 = p319 + tc;
                        p328 = p328 + tc;
                end
                335: begin
                        tc = f334;
                        p316 = p316 - tc;
                        p328 = p328 + tc;
                end
                336: begin
                        tc = f335;
                        p329 = p329 - tc;
                        p327 = p327 + tc;
                end
                337: begin
                        tc = f336;
                        p323 = p323 - tc;
                        p317 = p317 + tc;
                end
                338: begin
                        tc = f337;
                        p330 = p330 - tc;
                        p329 = p329 + tc;
                end
                339: begin
                        tc = f338;
                        p328 = p328 - tc;
                        p316 = p316 + tc*2;
                end
                340: begin
                        tc = f339;
                        p318 = p318 - tc;
                        p325 = p325 - tc;
                        p326 = p326 + tc;
                        p330 = p330 + tc;
                end
                341: begin
                        tc = f340;
                        p318 = p318 - tc;
                        p330 = p330 + tc;
                end
                342: begin
                        tc = f341;
                        p44 = p44 - tc;
                        p316 = p316 + tc;
                        p331 = p331 + tc;
                end
                343: begin
                        tc = f342;
                        p331 = p331 - tc;
                        p44 = p44 + tc;
                end
                344: begin
                        tc = f343;
                        p333 = p333 - tc;
                        p332 = p332 + tc;
                end
                345: begin
                        tc = f344;
                        p334 = p334 - tc;
                        p333 = p333 + tc;
                end
                346: begin
                        tc = f345;
                        p45 = p45 - tc;
                        p317 = p317 + tc;
                        p335 = p335 + tc;
                end
                347: begin
                        tc = f346;
                        p335 = p335 - tc;
                        p45 = p45 + tc;
                end
                348: begin
                        tc = f347;
                        p337 = p337 - tc;
                        p336 = p336 + tc;
                end
                349: begin
                        tc = f348;
                        p338 = p338 - tc;
                        p337 = p337 + tc;
                end
                350: begin
                        tc = f349;
                        p332 = p332 - tc;
                        p336 = p336 - tc;
                        p11 = p11 + tc;
                end
                351: begin
                        tc = f350;
                        p318 = p318 - tc;
                        p334 = p334 + tc;
                        p338 = p338 + tc;
                end
                352: begin
                        tc = f351;
                        p319 = p319 - tc;
                        p46 = p46 + tc;
                end
                353: begin
                        tc = f352;
                        p46 = p46 - tc;
                end
                354: begin
                        tc = f353;
                        p339 = p339 - tc;
                        p320 = p320 + tc;
                end
                355: begin
                        tc = f354;
                        p12 = p12 - tc;
                        p339 = p339 + tc;
                end
                356: begin
                        tc = f355;
                        p346 = p346 - tc;
                        p342 = p342 + tc;
                end
                357: begin
                        tc = f356;
                        p340 = p340 - tc;
                end
                358: begin
                        tc = f357;
                        p344 = p344 - tc;
                        p346 = p346 + tc;
                end
                359: begin
                        tc = f358;
                        p341 = p341 - tc*2;
                        p347 = p347 + tc;
                end
                360: begin
                        tc = f359;
                        p348 = p348 - tc;
                        p345 = p345 + tc;
                end
                361: begin
                        tc = f360;
                        p341 = p341 - tc;
                        p350 = p350 - tc;
                        p349 = p349 + tc;
                end
                362: begin
                        tc = f361;
                        p351 = p351 - tc;
                        p348 = p348 + tc;
                end
                363: begin
                        tc = f362;
                        p340 = p340 - tc;
                        p343 = p343 + tc;
                        p352 = p352 + tc;
                end
                364: begin
                        tc = f363;
                        p340 = p340 - tc;
                        p352 = p352 + tc;
                end
                365: begin
                        tc = f364;
                        p353 = p353 - tc;
                        p351 = p351 + tc;
                end
                366: begin
                        tc = f365;
                        p347 = p347 - tc;
                        p341 = p341 + tc;
                end
                367: begin
                        tc = f366;
                        p354 = p354 - tc;
                        p353 = p353 + tc;
                end
                368: begin
                        tc = f367;
                        p352 = p352 - tc;
                        p340 = p340 + tc*2;
                end
                369: begin
                        tc = f368;
                        p342 = p342 - tc;
                        p349 = p349 - tc;
                        p350 = p350 + tc;
                        p354 = p354 + tc;
                end
                370: begin
                        tc = f369;
                        p342 = p342 - tc;
                        p354 = p354 + tc;
                end
                371: begin
                        tc = f370;
                        p46 = p46 - tc;
                        p340 = p340 + tc;
                        p355 = p355 + tc;
                end
                372: begin
                        tc = f371;
                        p355 = p355 - tc;
                        p46 = p46 + tc;
                end
                373: begin
                        tc = f372;
                        p357 = p357 - tc;
                        p356 = p356 + tc;
                end
                374: begin
                        tc = f373;
                        p358 = p358 - tc;
                        p357 = p357 + tc;
                end
                375: begin
                        tc = f374;
                        p47 = p47 - tc;
                        p341 = p341 + tc;
                        p359 = p359 + tc;
                end
                376: begin
                        tc = f375;
                        p359 = p359 - tc;
                        p47 = p47 + tc;
                end
                377: begin
                        tc = f376;
                        p361 = p361 - tc;
                        p360 = p360 + tc;
                end
                378: begin
                        tc = f377;
                        p362 = p362 - tc;
                        p361 = p361 + tc;
                end
                379: begin
                        tc = f378;
                        p356 = p356 - tc;
                        p360 = p360 - tc;
                        p12 = p12 + tc;
                end
                380: begin
                        tc = f379;
                        p342 = p342 - tc;
                        p358 = p358 + tc;
                        p362 = p362 + tc;
                end
                381: begin
                        tc = f380;
                        p343 = p343 - tc;
                        p48 = p48 + tc;
                end
                382: begin
                        tc = f381;
                        p48 = p48 - tc;
                end
                383: begin
                        tc = f382;
                        p363 = p363 - tc;
                        p344 = p344 + tc;
                end
                384: begin
                        tc = f383;
                        p13 = p13 - tc;
                        p363 = p363 + tc;
                end
                385: begin
                        tc = f384;
                        p365 = p365 - tc;
                        p366 = p366 + tc;
                end
                386: begin
                        tc = f385;
                        p368 = p368 - tc;
                        p367 = p367 + tc;
                end
                387: begin
                        tc = f386;
                        p48 = p48 - tc;
                        p364 = p364 + tc;
                        p369 = p369 + tc;
                end
                388: begin
                        tc = f387;
                        p369 = p369 - tc;
                        p48 = p48 + tc;
                end
                389: begin
                        tc = f388;
                        p371 = p371 - tc;
                        p370 = p370 + tc;
                end
                390: begin
                        tc = f389;
                        p372 = p372 - tc;
                        p371 = p371 + tc;
                end
                391: begin
                        tc = f390;
                        p41 = p41 - tc;
                        p365 = p365 + tc;
                        p373 = p373 + tc;
                end
                392: begin
                        tc = f391;
                        p373 = p373 - tc;
                        p41 = p41 + tc;
                end
                393: begin
                        tc = f392;
                        p375 = p375 - tc;
                        p374 = p374 + tc;
                end
                394: begin
                        tc = f393;
                        p376 = p376 - tc;
                        p375 = p375 + tc;
                end
                395: begin
                        tc = f394;
                        p370 = p370 - tc;
                        p374 = p374 - tc;
                        p13 = p13 + tc;
                end
                396: begin
                        tc = f395;
                        p367 = p367 - tc;
                        p372 = p372 + tc;
                        p376 = p376 + tc;
                end
                397: begin
                        tc = f396;
                        p366 = p366 - tc;
                        p49 = p49 + tc;
                end
                398: begin
                        tc = f397;
                        p49 = p49 - tc;
                end
                399: begin
                        tc = f398;
                        p377 = p377 - tc;
                        p368 = p368 + tc;
                end
                400: begin
                        tc = f399;
                        p14 = p14 - tc;
                        p377 = p377 + tc;
                end
                401: begin
                        tc = f400;
                        p384 = p384 - tc;
                        p380 = p380 + tc;
                end
                402: begin
                        tc = f401;
                        p378 = p378 - tc;
                end
                403: begin
                        tc = f402;
                        p382 = p382 - tc;
                        p384 = p384 + tc;
                end
                404: begin
                        tc = f403;
                        p379 = p379 - tc*2;
                        p385 = p385 + tc;
                end
                405: begin
                        tc = f404;
                        p386 = p386 - tc;
                        p383 = p383 + tc;
                end
                406: begin
                        tc = f405;
                        p379 = p379 - tc;
                        p388 = p388 - tc;
                        p387 = p387 + tc;
                end
                407: begin
                        tc = f406;
                        p389 = p389 - tc;
                        p386 = p386 + tc;
                end
                408: begin
                        tc = f407;
                        p378 = p378 - tc;
                        p381 = p381 + tc;
                        p390 = p390 + tc;
                end
                409: begin
                        tc = f408;
                        p378 = p378 - tc;
                        p390 = p390 + tc;
                end
                410: begin
                        tc = f409;
                        p391 = p391 - tc;
                        p389 = p389 + tc;
                end
                411: begin
                        tc = f410;
                        p385 = p385 - tc;
                        p379 = p379 + tc;
                end
                412: begin
                        tc = f411;
                        p392 = p392 - tc;
                        p391 = p391 + tc;
                end
                413: begin
                        tc = f412;
                        p390 = p390 - tc;
                        p378 = p378 + tc*2;
                end
                414: begin
                        tc = f413;
                        p380 = p380 - tc;
                        p387 = p387 - tc;
                        p388 = p388 + tc;
                        p392 = p392 + tc;
                end
                415: begin
                        tc = f414;
                        p380 = p380 - tc;
                        p392 = p392 + tc;
                end
                416: begin
                        tc = f415;
                        p50 = p50 - tc;
                        p378 = p378 + tc;
                        p393 = p393 + tc;
                end
                417: begin
                        tc = f416;
                        p393 = p393 - tc;
                        p50 = p50 + tc;
                end
                418: begin
                        tc = f417;
                        p395 = p395 - tc;
                        p394 = p394 + tc;
                end
                419: begin
                        tc = f418;
                        p396 = p396 - tc;
                        p395 = p395 + tc;
                end
                420: begin
                        tc = f419;
                        p51 = p51 - tc;
                        p379 = p379 + tc;
                        p397 = p397 + tc;
                end
                421: begin
                        tc = f420;
                        p397 = p397 - tc;
                        p51 = p51 + tc;
                end
                422: begin
                        tc = f421;
                        p399 = p399 - tc;
                        p398 = p398 + tc;
                end
                423: begin
                        tc = f422;
                        p400 = p400 - tc;
                        p399 = p399 + tc;
                end
                424: begin
                        tc = f423;
                        p394 = p394 - tc;
                        p398 = p398 - tc;
                        p14 = p14 + tc;
                end
                425: begin
                        tc = f424;
                        p380 = p380 - tc;
                        p396 = p396 + tc;
                        p400 = p400 + tc;
                end
                426: begin
                        tc = f425;
                        p381 = p381 - tc;
                        p52 = p52 + tc;
                end
                427: begin
                        tc = f426;
                        p52 = p52 - tc;
                end
                428: begin
                        tc = f427;
                        p401 = p401 - tc;
                        p382 = p382 + tc;
                end
                429: begin
                        tc = f428;
                        p15 = p15 - tc;
                        p401 = p401 + tc;
                end
                430: begin
                        tc = f429;
                        p408 = p408 - tc;
                        p404 = p404 + tc;
                end
                431: begin
                        tc = f430;
                        p402 = p402 - tc;
                end
                432: begin
                        tc = f431;
                        p406 = p406 - tc;
                        p408 = p408 + tc;
                end
                433: begin
                        tc = f432;
                        p403 = p403 - tc*2;
                        p409 = p409 + tc;
                end
                434: begin
                        tc = f433;
                        p410 = p410 - tc;
                        p407 = p407 + tc;
                end
                435: begin
                        tc = f434;
                        p403 = p403 - tc;
                        p412 = p412 - tc;
                        p411 = p411 + tc;
                end
                436: begin
                        tc = f435;
                        p413 = p413 - tc;
                        p410 = p410 + tc;
                end
                437: begin
                        tc = f436;
                        p402 = p402 - tc;
                        p405 = p405 + tc;
                        p414 = p414 + tc;
                end
                438: begin
                        tc = f437;
                        p402 = p402 - tc;
                        p414 = p414 + tc;
                end
                439: begin
                        tc = f438;
                        p415 = p415 - tc;
                        p413 = p413 + tc;
                end
                440: begin
                        tc = f439;
                        p409 = p409 - tc;
                        p403 = p403 + tc;
                end
                441: begin
                        tc = f440;
                        p416 = p416 - tc;
                        p415 = p415 + tc;
                end
                442: begin
                        tc = f441;
                        p414 = p414 - tc;
                        p402 = p402 + tc*2;
                end
                443: begin
                        tc = f442;
                        p404 = p404 - tc;
                        p411 = p411 - tc;
                        p412 = p412 + tc;
                        p416 = p416 + tc;
                end
                444: begin
                        tc = f443;
                        p404 = p404 - tc;
                        p416 = p416 + tc;
                end
                445: begin
                        tc = f444;
                        p52 = p52 - tc;
                        p402 = p402 + tc;
                        p417 = p417 + tc;
                end
                446: begin
                        tc = f445;
                        p417 = p417 - tc;
                        p52 = p52 + tc;
                end
                447: begin
                        tc = f446;
                        p419 = p419 - tc;
                        p418 = p418 + tc;
                end
                448: begin
                        tc = f447;
                        p420 = p420 - tc;
                        p419 = p419 + tc;
                end
                449: begin
                        tc = f448;
                        p53 = p53 - tc;
                        p403 = p403 + tc;
                        p421 = p421 + tc;
                end
                450: begin
                        tc = f449;
                        p421 = p421 - tc;
                        p53 = p53 + tc;
                end
                451: begin
                        tc = f450;
                        p423 = p423 - tc;
                        p422 = p422 + tc;
                end
                452: begin
                        tc = f451;
                        p424 = p424 - tc;
                        p423 = p423 + tc;
                end
                453: begin
                        tc = f452;
                        p418 = p418 - tc;
                        p422 = p422 - tc;
                        p15 = p15 + tc;
                end
                454: begin
                        tc = f453;
                        p404 = p404 - tc;
                        p420 = p420 + tc;
                        p424 = p424 + tc;
                end
                455: begin
                        tc = f454;
                        p405 = p405 - tc;
                        p54 = p54 + tc;
                end
                456: begin
                        tc = f455;
                        p54 = p54 - tc;
                end
                457: begin
                        tc = f456;
                        p425 = p425 - tc;
                        p406 = p406 + tc;
                end
                458: begin
                        tc = f457;
                        p16 = p16 - tc;
                        p425 = p425 + tc;
                end
                459: begin
                        tc = f458;
                        p427 = p427 - tc;
                        p428 = p428 + tc;
                end
                460: begin
                        tc = f459;
                        p430 = p430 - tc;
                        p429 = p429 + tc;
                end
                461: begin
                        tc = f460;
                        p54 = p54 - tc;
                        p426 = p426 + tc;
                        p431 = p431 + tc;
                end
                462: begin
                        tc = f461;
                        p431 = p431 - tc;
                        p54 = p54 + tc;
                end
                463: begin
                        tc = f462;
                        p433 = p433 - tc;
                        p432 = p432 + tc;
                end
                464: begin
                        tc = f463;
                        p434 = p434 - tc;
                        p433 = p433 + tc;
                end
                465: begin
                        tc = f464;
                        p49 = p49 - tc;
                        p427 = p427 + tc;
                        p435 = p435 + tc;
                end
                466: begin
                        tc = f465;
                        p435 = p435 - tc;
                        p49 = p49 + tc;
                end
                467: begin
                        tc = f466;
                        p437 = p437 - tc;
                        p436 = p436 + tc;
                end
                468: begin
                        tc = f467;
                        p438 = p438 - tc;
                        p437 = p437 + tc;
                end
                469: begin
                        tc = f468;
                        p432 = p432 - tc;
                        p436 = p436 - tc;
                        p16 = p16 + tc;
                end
                470: begin
                        tc = f469;
                        p429 = p429 - tc;
                        p434 = p434 + tc;
                        p438 = p438 + tc;
                end
                471: begin
                        tc = f470;
                        p428 = p428 - tc;
                        p55 = p55 + tc;
                end
                472: begin
                        tc = f471;
                        p55 = p55 - tc;
                end
                473: begin
                        tc = f472;
                        p439 = p439 - tc;
                        p430 = p430 + tc;
                end
                474: begin
                        tc = f473;
                        p17 = p17 - tc;
                        p439 = p439 + tc;
                end
                475: begin
                        tc = f474;
                        p446 = p446 - tc;
                        p442 = p442 + tc;
                end
                476: begin
                        tc = f475;
                        p440 = p440 - tc;
                end
                477: begin
                        tc = f476;
                        p444 = p444 - tc;
                        p446 = p446 + tc;
                end
                478: begin
                        tc = f477;
                        p441 = p441 - tc*2;
                        p447 = p447 + tc;
                end
                479: begin
                        tc = f478;
                        p448 = p448 - tc;
                        p445 = p445 + tc;
                end
                480: begin
                        tc = f479;
                        p441 = p441 - tc;
                        p450 = p450 - tc;
                        p449 = p449 + tc;
                end
                481: begin
                        tc = f480;
                        p451 = p451 - tc;
                        p448 = p448 + tc;
                end
                482: begin
                        tc = f481;
                        p440 = p440 - tc;
                        p443 = p443 + tc;
                        p452 = p452 + tc;
                end
                483: begin
                        tc = f482;
                        p440 = p440 - tc;
                        p452 = p452 + tc;
                end
                484: begin
                        tc = f483;
                        p453 = p453 - tc;
                        p451 = p451 + tc;
                end
                485: begin
                        tc = f484;
                        p447 = p447 - tc;
                        p441 = p441 + tc;
                end
                486: begin
                        tc = f485;
                        p454 = p454 - tc;
                        p453 = p453 + tc;
                end
                487: begin
                        tc = f486;
                        p452 = p452 - tc;
                        p440 = p440 + tc*2;
                end
                488: begin
                        tc = f487;
                        p442 = p442 - tc;
                        p449 = p449 - tc;
                        p450 = p450 + tc;
                        p454 = p454 + tc;
                end
                489: begin
                        tc = f488;
                        p442 = p442 - tc;
                        p454 = p454 + tc;
                end
                490: begin
                        tc = f489;
                        p56 = p56 - tc;
                        p440 = p440 + tc;
                        p455 = p455 + tc;
                end
                491: begin
                        tc = f490;
                        p455 = p455 - tc;
                        p56 = p56 + tc;
                end
                492: begin
                        tc = f491;
                        p457 = p457 - tc;
                        p456 = p456 + tc;
                end
                493: begin
                        tc = f492;
                        p458 = p458 - tc;
                        p457 = p457 + tc;
                end
                494: begin
                        tc = f493;
                        p57 = p57 - tc;
                        p441 = p441 + tc;
                        p459 = p459 + tc;
                end
                495: begin
                        tc = f494;
                        p459 = p459 - tc;
                        p57 = p57 + tc;
                end
                496: begin
                        tc = f495;
                        p461 = p461 - tc;
                        p460 = p460 + tc;
                end
                497: begin
                        tc = f496;
                        p462 = p462 - tc;
                        p461 = p461 + tc;
                end
                498: begin
                        tc = f497;
                        p456 = p456 - tc;
                        p460 = p460 - tc;
                        p17 = p17 + tc;
                end
                499: begin
                        tc = f498;
                        p442 = p442 - tc;
                        p458 = p458 + tc;
                        p462 = p462 + tc;
                end
                500: begin
                        tc = f499;
                        p443 = p443 - tc;
                        p58 = p58 + tc;
                end
                501: begin
                        tc = f500;
                        p58 = p58 - tc;
                end
                502: begin
                        tc = f501;
                        p463 = p463 - tc;
                        p444 = p444 + tc;
                end
                503: begin
                        tc = f502;
                        p18 = p18 - tc;
                        p463 = p463 + tc;
                end
                504: begin
                        tc = f503;
                        p465 = p465 - tc;
                        p466 = p466 + tc;
                end
                505: begin
                        tc = f504;
                        p468 = p468 - tc;
                        p467 = p467 + tc;
                end
                506: begin
                        tc = f505;
                        p58 = p58 - tc;
                        p464 = p464 + tc;
                        p469 = p469 + tc;
                end
                507: begin
                        tc = f506;
                        p469 = p469 - tc;
                        p58 = p58 + tc;
                end
                508: begin
                        tc = f507;
                        p471 = p471 - tc;
                        p470 = p470 + tc;
                end
                509: begin
                        tc = f508;
                        p472 = p472 - tc;
                        p471 = p471 + tc;
                end
                510: begin
                        tc = f509;
                        p55 = p55 - tc;
                        p465 = p465 + tc;
                        p473 = p473 + tc;
                end
                511: begin
                        tc = f510;
                        p473 = p473 - tc;
                        p55 = p55 + tc;
                end
                512: begin
                        tc = f511;
                        p475 = p475 - tc;
                        p474 = p474 + tc;
                end
                513: begin
                        tc = f512;
                        p476 = p476 - tc;
                        p475 = p475 + tc;
                end
                514: begin
                        tc = f513;
                        p470 = p470 - tc;
                        p474 = p474 - tc;
                        p18 = p18 + tc;
                end
                515: begin
                        tc = f514;
                        p467 = p467 - tc;
                        p472 = p472 + tc;
                        p476 = p476 + tc;
                end
                516: begin
                        tc = f515;
                        p466 = p466 - tc;
                        p59 = p59 + tc;
                end
                517: begin
                        tc = f516;
                        p59 = p59 - tc;
                end
                518: begin
                        tc = f517;
                        p477 = p477 - tc;
                        p468 = p468 + tc;
                end
                519: begin
                        tc = f518;
                        p19 = p19 - tc;
                        p477 = p477 + tc;
                end
                520: begin
                        tc = f519;
                        p479 = p479 - tc;
                        p480 = p480 + tc;
                end
                521: begin
                        tc = f520;
                        p482 = p482 - tc;
                        p481 = p481 + tc;
                end
                522: begin
                        tc = f521;
                        p59 = p59 - tc;
                        p478 = p478 + tc;
                        p483 = p483 + tc;
                end
                523: begin
                        tc = f522;
                        p483 = p483 - tc;
                        p59 = p59 + tc;
                end
                524: begin
                        tc = f523;
                        p485 = p485 - tc;
                        p484 = p484 + tc;
                end
                525: begin
                        tc = f524;
                        p486 = p486 - tc;
                        p485 = p485 + tc;
                end
                526: begin
                        tc = f525;
                        p60 = p60 - tc;
                        p479 = p479 + tc;
                        p487 = p487 + tc;
                end
                527: begin
                        tc = f526;
                        p487 = p487 - tc;
                        p60 = p60 + tc;
                end
                528: begin
                        tc = f527;
                        p489 = p489 - tc;
                        p488 = p488 + tc;
                end
                529: begin
                        tc = f528;
                        p490 = p490 - tc;
                        p489 = p489 + tc;
                end
                530: begin
                        tc = f529;
                        p484 = p484 - tc;
                        p488 = p488 - tc;
                        p19 = p19 + tc;
                end
                531: begin
                        tc = f530;
                        p481 = p481 - tc;
                        p486 = p486 + tc;
                        p490 = p490 + tc;
                end
                532: begin
                        tc = f531;
                        p480 = p480 - tc;
                        p61 = p61 + tc;
                end
                533: begin
                        tc = f532;
                        p61 = p61 - tc;
                end
                534: begin
                        tc = f533;
                        p491 = p491 - tc;
                        p482 = p482 + tc;
                end
                535: begin
                        tc = f534;
                        p20 = p20 - tc;
                        p491 = p491 + tc;
                end
                default:;
        endcase
//        led = ~p61[9:6];
        if(tf>0) counter1=counter1+1;
end
end
reg [32:0] counter;

always @(posedge clk) begin
    if (counter < 32'd2_7500_0000)       //delay
        counter <= counter + 1'b1;
    else
        counter <= 32'd0;
end

always @(posedge clk) begin
    if (counter == 32'd0)       
        led <= ~counter1[47:42];
    else if (counter == 32'd2500_0000)       
        led <= ~counter1[41:36];
    else if (counter == 32'd5000_0000)       
        led <= ~counter1[35:30];
    else if (counter == 32'd7500_0000)       
        led <= ~counter1[29:24];
    else if (counter == 32'd1_0000_0000)       
        led <= ~counter1[23:18];
    else if (counter == 32'd1_2500_0000)       
        led <= ~counter1[17:12];
    else if (counter == 32'd1_5000_0000)       
        led <= ~counter1[11:6];
    else if (counter == 32'd1_7500_0000)       
        led <= ~counter1[5:0];
    else if (counter == 32'd2_0000_0000)       
        led <= 6'b000000;
    else if (counter == 32'd2_2500_0000)       
        led <= 6'b111111;
    else if (counter == 32'd2_5000_0000)       
        led <= 6'b000000;
    else
        led <= led;
end
endmodule