module sn(
        input clk,
        output reg [5:0] led
);
`define INH(place) ((place) == 0 ? 2047 : 0)
reg [10:0] p0=0,p1=1,p2=1,p3=1,p4=1,p5=1,p6=22,p7=33,p8=0,p9=25,p10=30,p11=0,p12=0,p13=1,p14=1,p15=1,p16=1,p17=22,p18=26,p19=0,p20=25,p21=34,p22=0,p23=0,p24=1,p25=1,p26=1,p27=1,p28=30,p29=33,p30=0,p31=29,p32=30,p33=0,p34=0,p35=1,p36=1,p37=1,p38=1,p39=30,p40=26,p41=0,p42=29,p43=34,p44=0,p45=0,p46=0,p47=0,p48=1,p49=0,p50=1,p51=1,p52=1,p53=0,p54=1,p55=0,p56=1,p57=1,p58=0,p59=1,p60=1,p61=0,p62=1,p63=1,p64=1,p65=0,p66=1,p67=1,p68=1,p69=1,p70=0,p71=0,p72=1,p73=0,p74=1,p75=1,p76=1,p77=0,p78=1,p79=0,p80=1,p81=1,p82=0,p83=1,p84=1,p85=0,p86=1,p87=1,p88=1,p89=0,p90=1,p91=1,p92=1,p93=1,p94=0,p95=0,p96=0,p97=1,p98=1,p99=0,p100=1,p101=1,p102=1,p103=0,p104=1,p105=1,p106=1,p107=1,p108=0,p109=0,p110=1,p111=0,p112=1,p113=1,p114=1,p115=0,p116=1,p117=0,p118=1,p119=1,p120=0,p121=1,p122=1,p123=0,p124=1,p125=1,p126=1,p127=0,p128=1,p129=1,p130=1,p131=1,p132=0,p133=0,p134=1,p135=0,p136=1,p137=1,p138=1,p139=0,p140=1,p141=0,p142=1,p143=1,p144=0,p145=1,p146=1,p147=0,p148=1,p149=1,p150=1,p151=0,p152=1,p153=1,p154=1,p155=1,p156=0,p157=0,p158=0,p159=1,p160=1,p161=0,p162=1,p163=1,p164=1,p165=0,p166=1,p167=1,p168=1,p169=1,p170=0,p171=0,p172=1,p173=0,p174=1,p175=1,p176=1,p177=0,p178=1,p179=0,p180=1,p181=1,p182=0,p183=1,p184=1,p185=0,p186=1,p187=1,p188=1,p189=0,p190=1,p191=1,p192=1,p193=1,p194=0,p195=0,p196=1,p197=0,p198=1,p199=1,p200=1,p201=0,p202=1,p203=0,p204=1,p205=1,p206=0,p207=1,p208=1,p209=0,p210=1,p211=1,p212=1,p213=0,p214=1,p215=1,p216=1,p217=1,p218=0,p219=0,p220=0,p221=1,p222=1,p223=0,p224=1,p225=1,p226=1,p227=0,p228=1,p229=1,p230=1,p231=1,p232=0,p233=0,p234=1,p235=0,p236=1,p237=1,p238=1,p239=0,p240=1,p241=0,p242=1,p243=1,p244=0,p245=1,p246=1,p247=0,p248=1,p249=1,p250=1,p251=0,p252=1,p253=1,p254=1,p255=1,p256=0,p257=0,p258=1,p259=0,p260=1,p261=1,p262=1,p263=0,p264=1,p265=0,p266=1,p267=1,p268=0,p269=1,p270=1,p271=0,p272=1,p273=1,p274=1,p275=0,p276=1,p277=1,p278=1,p279=1,p280=0,p281=0,p282=0,p283=1,p284=1,p285=0,p286=1,p287=1,p288=1,p289=0,p290=1,p291=1,p292=1,p293=1;
reg [10:0] f0,f1,f2,f3,f4,f5,f6,f7,f8,f9,f10,f11,f12,f13,f14,f15,f16,f17,f18,f19,f20,f21,f22,f23,f24,f25,f26,f27,f28,f29,f30,f31,f32,f33,f34,f35,f36,f37,f38,f39,f40,f41,f42,f43,f44,f45,f46,f47,f48,f49,f50,f51,f52,f53,f54,f55,f56,f57,f58,f59,f60,f61,f62,f63,f64,f65,f66,f67,f68,f69,f70,f71,f72,f73,f74,f75,f76,f77,f78,f79,f80,f81,f82,f83,f84,f85,f86,f87,f88,f89,f90,f91,f92,f93,f94,f95,f96,f97,f98,f99,f100,f101,f102,f103,f104,f105,f106,f107,f108,f109,f110,f111,f112,f113,f114,f115,f116,f117,f118,f119,f120,f121,f122,f123,f124,f125,f126,f127,f128,f129,f130,f131,f132,f133,f134,f135,f136,f137,f138,f139,f140,f141,f142,f143,f144,f145,f146,f147,f148,f149,f150,f151,f152,f153,f154,f155,f156,f157,f158,f159,f160,f161,f162,f163,f164,f165,f166,f167,f168,f169,f170,f171,f172,f173,f174,f175,f176,f177,f178,f179,f180,f181,f182,f183,f184,f185,f186,f187,f188,f189,f190,f191,f192,f193,f194,f195,f196,f197,f198,f199,f200,f201,f202,f203,f204,f205,f206,f207,f208,f209,f210,f211,f212,f213,f214,f215,f216,f217,f218,f219,f220,f221,f222,f223,f224,f225,f226,f227,f228,f229,f230,f231,f232,f233,f234,f235,f236,f237,f238,f239,f240,f241,f242,f243,f244,f245,f246,f247,f248,f249,f250,f251,f252,f253,f254,f255,f256,f257,f258,f259,f260,f261,f262,f263,f264,f265,f266,f267,f268,f269,f270,f271,f272,f273,f274,f275,f276,f277,f278,f279,f280,f281,f282,f283,f284,f285,f286,f287,f288,f289,f290,f291,f292,f293,f294,f295,f296,f297,f298,f299,f300,f301,f302,f303,f304,f305,f306,f307,f308,f309;
reg [10:0] tf;
reg [10:0] tc;
reg [1:0] clk_div; // 2位寄存器用于实现时钟分频
reg [47:0] counter1=1;
always @(posedge clk) begin
    if(clk_div < 2'b01)
        clk_div <= clk_div + 1; // 计数器自增
    else
        clk_div <= 2'b00; // 重置计数器
end

// 使用clk_div来控制某些逻辑的触发条件
always @(posedge clk) begin
    if (clk_div == 2'b01) begin
        f0 = 2047;
        f0 = (f0 >= `INH(p0)) ? `INH(p0) : f0;
        f0 = (f0 > p2) ? p2 : f0;
        f0 = (f0 > p13) ? p13 : f0;
        f0 = (f0 > p24) ? p24 : f0;
        f0 = (f0 > p35) ? p35 : f0;
        f1 = 2047;
        f1 = (f1 > p1) ? p1 : f1;
        f1 = (f1 >= `INH(p5)) ? `INH(p5) : f1;
        f1 = (f1 >= `INH(p16)) ? `INH(p16) : f1;
        f1 = (f1 >= `INH(p27)) ? `INH(p27) : f1;
        f1 = (f1 >= `INH(p38)) ? `INH(p38) : f1;
        f2 = 2047;
        f2 = (f2 >= `INH(p48)) ? `INH(p48) : f2;
        f2 = (f2 > p51) ? p51 : f2;
        f3 = 2047;
        f3 = (f3 >= `INH(p72)) ? `INH(p72) : f3;
        f3 = (f3 > p75) ? p75 : f3;
        f4 = 2047;
        f4 = (f4 > p94) ? p94 : f4;
        f4 = (f4 >= `INH(p97)) ? `INH(p97) : f4;
        f5 = 2047;
        f5 = (f5 >= `INH(p110)) ? `INH(p110) : f5;
        f5 = (f5 > p113) ? p113 : f5;
        f6 = 2047;
        f6 = (f6 >= `INH(p134)) ? `INH(p134) : f6;
        f6 = (f6 > p137) ? p137 : f6;
        f7 = 2047;
        f7 = (f7 > p156) ? p156 : f7;
        f7 = (f7 >= `INH(p159)) ? `INH(p159) : f7;
        f8 = 2047;
        f8 = (f8 >= `INH(p172)) ? `INH(p172) : f8;
        f8 = (f8 > p175) ? p175 : f8;
        f9 = 2047;
        f9 = (f9 >= `INH(p196)) ? `INH(p196) : f9;
        f9 = (f9 > p199) ? p199 : f9;
        f10 = 2047;
        f10 = (f10 > p218) ? p218 : f10;
        f10 = (f10 >= `INH(p221)) ? `INH(p221) : f10;
        f11 = 2047;
        f11 = (f11 >= `INH(p234)) ? `INH(p234) : f11;
        f11 = (f11 > p237) ? p237 : f11;
        f12 = 2047;
        f12 = (f12 >= `INH(p258)) ? `INH(p258) : f12;
        f12 = (f12 > p261) ? p261 : f12;
        f13 = 2047;
        f13 = (f13 > p280) ? p280 : f13;
        f13 = (f13 >= `INH(p283)) ? `INH(p283) : f13;
        f14 = 2047;
        f14 = (f14 >= `INH(p47)) ? `INH(p47) : f14;
        f14 = (f14 >= `INH(p48)) ? `INH(p48) : f14;
        f14 = (f14 > p52) ? p52 : f14;
        f15 = 2047;
        f15 = (f15 > p46) ? p46 : f15;
        f15 = (f15 >= `INH(p52)) ? `INH(p52) : f15;
        f16 = 2047;
        f16 = (f16 > p50) ? p50 : f16;
        f16 = (f16 >= `INH(p52)) ? `INH(p52) : f16;
        f17 = 2047;
        f17 = (f17 >= p47/2) ? p47/2 : f17;
        f17 = (f17 >= `INH(p51)) ? `INH(p51) : f17;
        f18 = 2047;
        f18 = (f18 >= `INH(p51)) ? `INH(p51) : f18;
        f18 = (f18 > p54) ? p54 : f18;
        f19 = 2047;
        f19 = (f19 > p47) ? p47 : f19;
        f19 = (f19 >= `INH(p54)) ? `INH(p54) : f19;
        f19 = (f19 > p56) ? p56 : f19;
        f20 = 2047;
        f20 = (f20 >= `INH(p54)) ? `INH(p54) : f20;
        f20 = (f20 > p57) ? p57 : f20;
        f21 = 2047;
        f21 = (f21 > p46) ? p46 : f21;
        f21 = (f21 >= `INH(p56)) ? `INH(p56) : f21;
        f21 = (f21 >= `INH(p57)) ? `INH(p57) : f21;
        f22 = 2047;
        f22 = (f22 > p46) ? p46 : f22;
        f22 = (f22 >= `INH(p55)) ? `INH(p55) : f22;
        f22 = (f22 >= `INH(p57)) ? `INH(p57) : f22;
        f23 = 2047;
        f23 = (f23 >= `INH(p57)) ? `INH(p57) : f23;
        f23 = (f23 > p59) ? p59 : f23;
        f24 = 2047;
        f24 = (f24 > p53) ? p53 : f24;
        f24 = (f24 >= `INH(p59)) ? `INH(p59) : f24;
        f25 = 2047;
        f25 = (f25 >= `INH(p59)) ? `INH(p59) : f25;
        f25 = (f25 > p60) ? p60 : f25;
        f26 = 2047;
        f26 = (f26 > p58) ? p58 : f26;
        f26 = (f26 >= `INH(p60)) ? `INH(p60) : f26;
        f27 = 2047;
        f27 = (f27 > p48) ? p48 : f27;
        f27 = (f27 > p55) ? p55 : f27;
        f27 = (f27 >= `INH(p56)) ? `INH(p56) : f27;
        f27 = (f27 >= `INH(p60)) ? `INH(p60) : f27;
        f28 = 2047;
        f28 = (f28 > p48) ? p48 : f28;
        f28 = (f28 >= `INH(p55)) ? `INH(p55) : f28;
        f28 = (f28 >= `INH(p60)) ? `INH(p60) : f28;
        f29 = 2047;
        f29 = (f29 > p6) ? p6 : f29;
        f29 = (f29 >= `INH(p62)) ? `INH(p62) : f29;
        f30 = 2047;
        f30 = (f30 > p61) ? p61 : f30;
        f30 = (f30 >= `INH(p63)) ? `INH(p63) : f30;
        f31 = 2047;
        f31 = (f31 >= `INH(p6)) ? `INH(p6) : f31;
        f31 = (f31 >= `INH(p62)) ? `INH(p62) : f31;
        f31 = (f31 > p63) ? p63 : f31;
        f32 = 2047;
        f32 = (f32 >= `INH(p61)) ? `INH(p61) : f32;
        f32 = (f32 >= `INH(p63)) ? `INH(p63) : f32;
        f32 = (f32 > p64) ? p64 : f32;
        f33 = 2047;
        f33 = (f33 > p7) ? p7 : f33;
        f33 = (f33 >= `INH(p66)) ? `INH(p66) : f33;
        f34 = 2047;
        f34 = (f34 > p65) ? p65 : f34;
        f34 = (f34 >= `INH(p67)) ? `INH(p67) : f34;
        f35 = 2047;
        f35 = (f35 >= `INH(p7)) ? `INH(p7) : f35;
        f35 = (f35 >= `INH(p66)) ? `INH(p66) : f35;
        f35 = (f35 > p67) ? p67 : f35;
        f36 = 2047;
        f36 = (f36 >= `INH(p65)) ? `INH(p65) : f36;
        f36 = (f36 >= `INH(p67)) ? `INH(p67) : f36;
        f36 = (f36 > p68) ? p68 : f36;
        f37 = 2047;
        f37 = (f37 >= `INH(p2)) ? `INH(p2) : f37;
        f37 = (f37 > p62) ? p62 : f37;
        f37 = (f37 > p66) ? p66 : f37;
        f38 = 2047;
        f38 = (f38 > p48) ? p48 : f38;
        f38 = (f38 >= `INH(p64)) ? `INH(p64) : f38;
        f38 = (f38 >= `INH(p68)) ? `INH(p68) : f38;
        f39 = 2047;
        f39 = (f39 > p49) ? p49 : f39;
        f39 = (f39 >= `INH(p69)) ? `INH(p69) : f39;
        f40 = 2047;
        f40 = (f40 > p8) ? p8 : f40;
        f40 = (f40 >= `INH(p50)) ? `INH(p50) : f40;
        f41 = 2047;
        f41 = (f41 >= `INH(p8)) ? `INH(p8) : f41;
        f41 = (f41 >= `INH(p50)) ? `INH(p50) : f41;
        f41 = (f41 > p69) ? p69 : f41;
        f42 = 2047;
        f42 = (f42 > p3) ? p3 : f42;
        f42 = (f42 >= `INH(p49)) ? `INH(p49) : f42;
        f42 = (f42 >= `INH(p69)) ? `INH(p69) : f42;
        f43 = 2047;
        f43 = (f43 >= `INH(p71)) ? `INH(p71) : f43;
        f43 = (f43 >= `INH(p72)) ? `INH(p72) : f43;
        f43 = (f43 > p76) ? p76 : f43;
        f44 = 2047;
        f44 = (f44 > p70) ? p70 : f44;
        f44 = (f44 >= `INH(p76)) ? `INH(p76) : f44;
        f45 = 2047;
        f45 = (f45 > p74) ? p74 : f45;
        f45 = (f45 >= `INH(p76)) ? `INH(p76) : f45;
        f46 = 2047;
        f46 = (f46 >= p71/2) ? p71/2 : f46;
        f46 = (f46 >= `INH(p75)) ? `INH(p75) : f46;
        f47 = 2047;
        f47 = (f47 >= `INH(p75)) ? `INH(p75) : f47;
        f47 = (f47 > p78) ? p78 : f47;
        f48 = 2047;
        f48 = (f48 > p71) ? p71 : f48;
        f48 = (f48 >= `INH(p78)) ? `INH(p78) : f48;
        f48 = (f48 > p80) ? p80 : f48;
        f49 = 2047;
        f49 = (f49 >= `INH(p78)) ? `INH(p78) : f49;
        f49 = (f49 > p81) ? p81 : f49;
        f50 = 2047;
        f50 = (f50 > p70) ? p70 : f50;
        f50 = (f50 >= `INH(p80)) ? `INH(p80) : f50;
        f50 = (f50 >= `INH(p81)) ? `INH(p81) : f50;
        f51 = 2047;
        f51 = (f51 > p70) ? p70 : f51;
        f51 = (f51 >= `INH(p79)) ? `INH(p79) : f51;
        f51 = (f51 >= `INH(p81)) ? `INH(p81) : f51;
        f52 = 2047;
        f52 = (f52 >= `INH(p81)) ? `INH(p81) : f52;
        f52 = (f52 > p83) ? p83 : f52;
        f53 = 2047;
        f53 = (f53 > p77) ? p77 : f53;
        f53 = (f53 >= `INH(p83)) ? `INH(p83) : f53;
        f54 = 2047;
        f54 = (f54 >= `INH(p83)) ? `INH(p83) : f54;
        f54 = (f54 > p84) ? p84 : f54;
        f55 = 2047;
        f55 = (f55 > p82) ? p82 : f55;
        f55 = (f55 >= `INH(p84)) ? `INH(p84) : f55;
        f56 = 2047;
        f56 = (f56 > p72) ? p72 : f56;
        f56 = (f56 > p79) ? p79 : f56;
        f56 = (f56 >= `INH(p80)) ? `INH(p80) : f56;
        f56 = (f56 >= `INH(p84)) ? `INH(p84) : f56;
        f57 = 2047;
        f57 = (f57 > p72) ? p72 : f57;
        f57 = (f57 >= `INH(p79)) ? `INH(p79) : f57;
        f57 = (f57 >= `INH(p84)) ? `INH(p84) : f57;
        f58 = 2047;
        f58 = (f58 > p9) ? p9 : f58;
        f58 = (f58 >= `INH(p86)) ? `INH(p86) : f58;
        f59 = 2047;
        f59 = (f59 > p85) ? p85 : f59;
        f59 = (f59 >= `INH(p87)) ? `INH(p87) : f59;
        f60 = 2047;
        f60 = (f60 >= `INH(p9)) ? `INH(p9) : f60;
        f60 = (f60 >= `INH(p86)) ? `INH(p86) : f60;
        f60 = (f60 > p87) ? p87 : f60;
        f61 = 2047;
        f61 = (f61 >= `INH(p85)) ? `INH(p85) : f61;
        f61 = (f61 >= `INH(p87)) ? `INH(p87) : f61;
        f61 = (f61 > p88) ? p88 : f61;
        f62 = 2047;
        f62 = (f62 > p10) ? p10 : f62;
        f62 = (f62 >= `INH(p90)) ? `INH(p90) : f62;
        f63 = 2047;
        f63 = (f63 > p89) ? p89 : f63;
        f63 = (f63 >= `INH(p91)) ? `INH(p91) : f63;
        f64 = 2047;
        f64 = (f64 >= `INH(p10)) ? `INH(p10) : f64;
        f64 = (f64 >= `INH(p90)) ? `INH(p90) : f64;
        f64 = (f64 > p91) ? p91 : f64;
        f65 = 2047;
        f65 = (f65 >= `INH(p89)) ? `INH(p89) : f65;
        f65 = (f65 >= `INH(p91)) ? `INH(p91) : f65;
        f65 = (f65 > p92) ? p92 : f65;
        f66 = 2047;
        f66 = (f66 >= `INH(p3)) ? `INH(p3) : f66;
        f66 = (f66 > p86) ? p86 : f66;
        f66 = (f66 > p90) ? p90 : f66;
        f67 = 2047;
        f67 = (f67 > p72) ? p72 : f67;
        f67 = (f67 >= `INH(p88)) ? `INH(p88) : f67;
        f67 = (f67 >= `INH(p92)) ? `INH(p92) : f67;
        f68 = 2047;
        f68 = (f68 > p73) ? p73 : f68;
        f68 = (f68 >= `INH(p93)) ? `INH(p93) : f68;
        f69 = 2047;
        f69 = (f69 > p11) ? p11 : f69;
        f69 = (f69 >= `INH(p74)) ? `INH(p74) : f69;
        f70 = 2047;
        f70 = (f70 >= `INH(p11)) ? `INH(p11) : f70;
        f70 = (f70 >= `INH(p74)) ? `INH(p74) : f70;
        f70 = (f70 > p93) ? p93 : f70;
        f71 = 2047;
        f71 = (f71 > p4) ? p4 : f71;
        f71 = (f71 >= `INH(p73)) ? `INH(p73) : f71;
        f71 = (f71 >= `INH(p93)) ? `INH(p93) : f71;
        f72 = 2047;
        f72 = (f72 > p95) ? p95 : f72;
        f72 = (f72 >= `INH(p97)) ? `INH(p97) : f72;
        f73 = 2047;
        f73 = (f73 >= `INH(p94)) ? `INH(p94) : f73;
        f73 = (f73 >= `INH(p95)) ? `INH(p95) : f73;
        f73 = (f73 >= `INH(p97)) ? `INH(p97) : f73;
        f73 = (f73 > p98) ? p98 : f73;
        f74 = 2047;
        f74 = (f74 > p8) ? p8 : f74;
        f74 = (f74 >= `INH(p100)) ? `INH(p100) : f74;
        f75 = 2047;
        f75 = (f75 > p99) ? p99 : f75;
        f75 = (f75 >= `INH(p101)) ? `INH(p101) : f75;
        f76 = 2047;
        f76 = (f76 >= `INH(p8)) ? `INH(p8) : f76;
        f76 = (f76 >= `INH(p100)) ? `INH(p100) : f76;
        f76 = (f76 > p101) ? p101 : f76;
        f77 = 2047;
        f77 = (f77 >= `INH(p99)) ? `INH(p99) : f77;
        f77 = (f77 >= `INH(p101)) ? `INH(p101) : f77;
        f77 = (f77 > p102) ? p102 : f77;
        f78 = 2047;
        f78 = (f78 > p11) ? p11 : f78;
        f78 = (f78 >= `INH(p104)) ? `INH(p104) : f78;
        f79 = 2047;
        f79 = (f79 > p103) ? p103 : f79;
        f79 = (f79 >= `INH(p105)) ? `INH(p105) : f79;
        f80 = 2047;
        f80 = (f80 >= `INH(p11)) ? `INH(p11) : f80;
        f80 = (f80 >= `INH(p104)) ? `INH(p104) : f80;
        f80 = (f80 > p105) ? p105 : f80;
        f81 = 2047;
        f81 = (f81 >= `INH(p103)) ? `INH(p103) : f81;
        f81 = (f81 >= `INH(p105)) ? `INH(p105) : f81;
        f81 = (f81 > p106) ? p106 : f81;
        f82 = 2047;
        f82 = (f82 >= `INH(p4)) ? `INH(p4) : f82;
        f82 = (f82 > p100) ? p100 : f82;
        f82 = (f82 > p104) ? p104 : f82;
        f83 = 2047;
        f83 = (f83 > p97) ? p97 : f83;
        f83 = (f83 >= `INH(p102)) ? `INH(p102) : f83;
        f83 = (f83 >= `INH(p106)) ? `INH(p106) : f83;
        f84 = 2047;
        f84 = (f84 > p96) ? p96 : f84;
        f84 = (f84 >= `INH(p107)) ? `INH(p107) : f84;
        f85 = 2047;
        f85 = (f85 > p12) ? p12 : f85;
        f85 = (f85 >= `INH(p98)) ? `INH(p98) : f85;
        f86 = 2047;
        f86 = (f86 >= `INH(p12)) ? `INH(p12) : f86;
        f86 = (f86 >= `INH(p98)) ? `INH(p98) : f86;
        f86 = (f86 > p107) ? p107 : f86;
        f87 = 2047;
        f87 = (f87 > p5) ? p5 : f87;
        f87 = (f87 >= `INH(p96)) ? `INH(p96) : f87;
        f87 = (f87 >= `INH(p107)) ? `INH(p107) : f87;
        f88 = 2047;
        f88 = (f88 >= `INH(p109)) ? `INH(p109) : f88;
        f88 = (f88 >= `INH(p110)) ? `INH(p110) : f88;
        f88 = (f88 > p114) ? p114 : f88;
        f89 = 2047;
        f89 = (f89 > p108) ? p108 : f89;
        f89 = (f89 >= `INH(p114)) ? `INH(p114) : f89;
        f90 = 2047;
        f90 = (f90 > p112) ? p112 : f90;
        f90 = (f90 >= `INH(p114)) ? `INH(p114) : f90;
        f91 = 2047;
        f91 = (f91 >= p109/2) ? p109/2 : f91;
        f91 = (f91 >= `INH(p113)) ? `INH(p113) : f91;
        f92 = 2047;
        f92 = (f92 >= `INH(p113)) ? `INH(p113) : f92;
        f92 = (f92 > p116) ? p116 : f92;
        f93 = 2047;
        f93 = (f93 > p109) ? p109 : f93;
        f93 = (f93 >= `INH(p116)) ? `INH(p116) : f93;
        f93 = (f93 > p118) ? p118 : f93;
        f94 = 2047;
        f94 = (f94 >= `INH(p116)) ? `INH(p116) : f94;
        f94 = (f94 > p119) ? p119 : f94;
        f95 = 2047;
        f95 = (f95 > p108) ? p108 : f95;
        f95 = (f95 >= `INH(p118)) ? `INH(p118) : f95;
        f95 = (f95 >= `INH(p119)) ? `INH(p119) : f95;
        f96 = 2047;
        f96 = (f96 > p108) ? p108 : f96;
        f96 = (f96 >= `INH(p117)) ? `INH(p117) : f96;
        f96 = (f96 >= `INH(p119)) ? `INH(p119) : f96;
        f97 = 2047;
        f97 = (f97 >= `INH(p119)) ? `INH(p119) : f97;
        f97 = (f97 > p121) ? p121 : f97;
        f98 = 2047;
        f98 = (f98 > p115) ? p115 : f98;
        f98 = (f98 >= `INH(p121)) ? `INH(p121) : f98;
        f99 = 2047;
        f99 = (f99 >= `INH(p121)) ? `INH(p121) : f99;
        f99 = (f99 > p122) ? p122 : f99;
        f100 = 2047;
        f100 = (f100 > p120) ? p120 : f100;
        f100 = (f100 >= `INH(p122)) ? `INH(p122) : f100;
        f101 = 2047;
        f101 = (f101 > p110) ? p110 : f101;
        f101 = (f101 > p117) ? p117 : f101;
        f101 = (f101 >= `INH(p118)) ? `INH(p118) : f101;
        f101 = (f101 >= `INH(p122)) ? `INH(p122) : f101;
        f102 = 2047;
        f102 = (f102 > p110) ? p110 : f102;
        f102 = (f102 >= `INH(p117)) ? `INH(p117) : f102;
        f102 = (f102 >= `INH(p122)) ? `INH(p122) : f102;
        f103 = 2047;
        f103 = (f103 > p17) ? p17 : f103;
        f103 = (f103 >= `INH(p124)) ? `INH(p124) : f103;
        f104 = 2047;
        f104 = (f104 > p123) ? p123 : f104;
        f104 = (f104 >= `INH(p125)) ? `INH(p125) : f104;
        f105 = 2047;
        f105 = (f105 >= `INH(p17)) ? `INH(p17) : f105;
        f105 = (f105 >= `INH(p124)) ? `INH(p124) : f105;
        f105 = (f105 > p125) ? p125 : f105;
        f106 = 2047;
        f106 = (f106 >= `INH(p123)) ? `INH(p123) : f106;
        f106 = (f106 >= `INH(p125)) ? `INH(p125) : f106;
        f106 = (f106 > p126) ? p126 : f106;
        f107 = 2047;
        f107 = (f107 > p18) ? p18 : f107;
        f107 = (f107 >= `INH(p128)) ? `INH(p128) : f107;
        f108 = 2047;
        f108 = (f108 > p127) ? p127 : f108;
        f108 = (f108 >= `INH(p129)) ? `INH(p129) : f108;
        f109 = 2047;
        f109 = (f109 >= `INH(p18)) ? `INH(p18) : f109;
        f109 = (f109 >= `INH(p128)) ? `INH(p128) : f109;
        f109 = (f109 > p129) ? p129 : f109;
        f110 = 2047;
        f110 = (f110 >= `INH(p127)) ? `INH(p127) : f110;
        f110 = (f110 >= `INH(p129)) ? `INH(p129) : f110;
        f110 = (f110 > p130) ? p130 : f110;
        f111 = 2047;
        f111 = (f111 >= `INH(p13)) ? `INH(p13) : f111;
        f111 = (f111 > p124) ? p124 : f111;
        f111 = (f111 > p128) ? p128 : f111;
        f112 = 2047;
        f112 = (f112 > p110) ? p110 : f112;
        f112 = (f112 >= `INH(p126)) ? `INH(p126) : f112;
        f112 = (f112 >= `INH(p130)) ? `INH(p130) : f112;
        f113 = 2047;
        f113 = (f113 > p111) ? p111 : f113;
        f113 = (f113 >= `INH(p131)) ? `INH(p131) : f113;
        f114 = 2047;
        f114 = (f114 > p19) ? p19 : f114;
        f114 = (f114 >= `INH(p112)) ? `INH(p112) : f114;
        f115 = 2047;
        f115 = (f115 >= `INH(p19)) ? `INH(p19) : f115;
        f115 = (f115 >= `INH(p112)) ? `INH(p112) : f115;
        f115 = (f115 > p131) ? p131 : f115;
        f116 = 2047;
        f116 = (f116 > p14) ? p14 : f116;
        f116 = (f116 >= `INH(p111)) ? `INH(p111) : f116;
        f116 = (f116 >= `INH(p131)) ? `INH(p131) : f116;
        f117 = 2047;
        f117 = (f117 >= `INH(p133)) ? `INH(p133) : f117;
        f117 = (f117 >= `INH(p134)) ? `INH(p134) : f117;
        f117 = (f117 > p138) ? p138 : f117;
        f118 = 2047;
        f118 = (f118 > p132) ? p132 : f118;
        f118 = (f118 >= `INH(p138)) ? `INH(p138) : f118;
        f119 = 2047;
        f119 = (f119 > p136) ? p136 : f119;
        f119 = (f119 >= `INH(p138)) ? `INH(p138) : f119;
        f120 = 2047;
        f120 = (f120 >= p133/2) ? p133/2 : f120;
        f120 = (f120 >= `INH(p137)) ? `INH(p137) : f120;
        f121 = 2047;
        f121 = (f121 >= `INH(p137)) ? `INH(p137) : f121;
        f121 = (f121 > p140) ? p140 : f121;
        f122 = 2047;
        f122 = (f122 > p133) ? p133 : f122;
        f122 = (f122 >= `INH(p140)) ? `INH(p140) : f122;
        f122 = (f122 > p142) ? p142 : f122;
        f123 = 2047;
        f123 = (f123 >= `INH(p140)) ? `INH(p140) : f123;
        f123 = (f123 > p143) ? p143 : f123;
        f124 = 2047;
        f124 = (f124 > p132) ? p132 : f124;
        f124 = (f124 >= `INH(p142)) ? `INH(p142) : f124;
        f124 = (f124 >= `INH(p143)) ? `INH(p143) : f124;
        f125 = 2047;
        f125 = (f125 > p132) ? p132 : f125;
        f125 = (f125 >= `INH(p141)) ? `INH(p141) : f125;
        f125 = (f125 >= `INH(p143)) ? `INH(p143) : f125;
        f126 = 2047;
        f126 = (f126 >= `INH(p143)) ? `INH(p143) : f126;
        f126 = (f126 > p145) ? p145 : f126;
        f127 = 2047;
        f127 = (f127 > p139) ? p139 : f127;
        f127 = (f127 >= `INH(p145)) ? `INH(p145) : f127;
        f128 = 2047;
        f128 = (f128 >= `INH(p145)) ? `INH(p145) : f128;
        f128 = (f128 > p146) ? p146 : f128;
        f129 = 2047;
        f129 = (f129 > p144) ? p144 : f129;
        f129 = (f129 >= `INH(p146)) ? `INH(p146) : f129;
        f130 = 2047;
        f130 = (f130 > p134) ? p134 : f130;
        f130 = (f130 > p141) ? p141 : f130;
        f130 = (f130 >= `INH(p142)) ? `INH(p142) : f130;
        f130 = (f130 >= `INH(p146)) ? `INH(p146) : f130;
        f131 = 2047;
        f131 = (f131 > p134) ? p134 : f131;
        f131 = (f131 >= `INH(p141)) ? `INH(p141) : f131;
        f131 = (f131 >= `INH(p146)) ? `INH(p146) : f131;
        f132 = 2047;
        f132 = (f132 > p20) ? p20 : f132;
        f132 = (f132 >= `INH(p148)) ? `INH(p148) : f132;
        f133 = 2047;
        f133 = (f133 > p147) ? p147 : f133;
        f133 = (f133 >= `INH(p149)) ? `INH(p149) : f133;
        f134 = 2047;
        f134 = (f134 >= `INH(p20)) ? `INH(p20) : f134;
        f134 = (f134 >= `INH(p148)) ? `INH(p148) : f134;
        f134 = (f134 > p149) ? p149 : f134;
        f135 = 2047;
        f135 = (f135 >= `INH(p147)) ? `INH(p147) : f135;
        f135 = (f135 >= `INH(p149)) ? `INH(p149) : f135;
        f135 = (f135 > p150) ? p150 : f135;
        f136 = 2047;
        f136 = (f136 > p21) ? p21 : f136;
        f136 = (f136 >= `INH(p152)) ? `INH(p152) : f136;
        f137 = 2047;
        f137 = (f137 > p151) ? p151 : f137;
        f137 = (f137 >= `INH(p153)) ? `INH(p153) : f137;
        f138 = 2047;
        f138 = (f138 >= `INH(p21)) ? `INH(p21) : f138;
        f138 = (f138 >= `INH(p152)) ? `INH(p152) : f138;
        f138 = (f138 > p153) ? p153 : f138;
        f139 = 2047;
        f139 = (f139 >= `INH(p151)) ? `INH(p151) : f139;
        f139 = (f139 >= `INH(p153)) ? `INH(p153) : f139;
        f139 = (f139 > p154) ? p154 : f139;
        f140 = 2047;
        f140 = (f140 >= `INH(p14)) ? `INH(p14) : f140;
        f140 = (f140 > p148) ? p148 : f140;
        f140 = (f140 > p152) ? p152 : f140;
        f141 = 2047;
        f141 = (f141 > p134) ? p134 : f141;
        f141 = (f141 >= `INH(p150)) ? `INH(p150) : f141;
        f141 = (f141 >= `INH(p154)) ? `INH(p154) : f141;
        f142 = 2047;
        f142 = (f142 > p135) ? p135 : f142;
        f142 = (f142 >= `INH(p155)) ? `INH(p155) : f142;
        f143 = 2047;
        f143 = (f143 > p22) ? p22 : f143;
        f143 = (f143 >= `INH(p136)) ? `INH(p136) : f143;
        f144 = 2047;
        f144 = (f144 >= `INH(p22)) ? `INH(p22) : f144;
        f144 = (f144 >= `INH(p136)) ? `INH(p136) : f144;
        f144 = (f144 > p155) ? p155 : f144;
        f145 = 2047;
        f145 = (f145 > p15) ? p15 : f145;
        f145 = (f145 >= `INH(p135)) ? `INH(p135) : f145;
        f145 = (f145 >= `INH(p155)) ? `INH(p155) : f145;
        f146 = 2047;
        f146 = (f146 > p157) ? p157 : f146;
        f146 = (f146 >= `INH(p159)) ? `INH(p159) : f146;
        f147 = 2047;
        f147 = (f147 >= `INH(p156)) ? `INH(p156) : f147;
        f147 = (f147 >= `INH(p157)) ? `INH(p157) : f147;
        f147 = (f147 >= `INH(p159)) ? `INH(p159) : f147;
        f147 = (f147 > p160) ? p160 : f147;
        f148 = 2047;
        f148 = (f148 > p19) ? p19 : f148;
        f148 = (f148 >= `INH(p162)) ? `INH(p162) : f148;
        f149 = 2047;
        f149 = (f149 > p161) ? p161 : f149;
        f149 = (f149 >= `INH(p163)) ? `INH(p163) : f149;
        f150 = 2047;
        f150 = (f150 >= `INH(p19)) ? `INH(p19) : f150;
        f150 = (f150 >= `INH(p162)) ? `INH(p162) : f150;
        f150 = (f150 > p163) ? p163 : f150;
        f151 = 2047;
        f151 = (f151 >= `INH(p161)) ? `INH(p161) : f151;
        f151 = (f151 >= `INH(p163)) ? `INH(p163) : f151;
        f151 = (f151 > p164) ? p164 : f151;
        f152 = 2047;
        f152 = (f152 > p22) ? p22 : f152;
        f152 = (f152 >= `INH(p166)) ? `INH(p166) : f152;
        f153 = 2047;
        f153 = (f153 > p165) ? p165 : f153;
        f153 = (f153 >= `INH(p167)) ? `INH(p167) : f153;
        f154 = 2047;
        f154 = (f154 >= `INH(p22)) ? `INH(p22) : f154;
        f154 = (f154 >= `INH(p166)) ? `INH(p166) : f154;
        f154 = (f154 > p167) ? p167 : f154;
        f155 = 2047;
        f155 = (f155 >= `INH(p165)) ? `INH(p165) : f155;
        f155 = (f155 >= `INH(p167)) ? `INH(p167) : f155;
        f155 = (f155 > p168) ? p168 : f155;
        f156 = 2047;
        f156 = (f156 >= `INH(p15)) ? `INH(p15) : f156;
        f156 = (f156 > p162) ? p162 : f156;
        f156 = (f156 > p166) ? p166 : f156;
        f157 = 2047;
        f157 = (f157 > p159) ? p159 : f157;
        f157 = (f157 >= `INH(p164)) ? `INH(p164) : f157;
        f157 = (f157 >= `INH(p168)) ? `INH(p168) : f157;
        f158 = 2047;
        f158 = (f158 > p158) ? p158 : f158;
        f158 = (f158 >= `INH(p169)) ? `INH(p169) : f158;
        f159 = 2047;
        f159 = (f159 > p23) ? p23 : f159;
        f159 = (f159 >= `INH(p160)) ? `INH(p160) : f159;
        f160 = 2047;
        f160 = (f160 >= `INH(p23)) ? `INH(p23) : f160;
        f160 = (f160 >= `INH(p160)) ? `INH(p160) : f160;
        f160 = (f160 > p169) ? p169 : f160;
        f161 = 2047;
        f161 = (f161 > p16) ? p16 : f161;
        f161 = (f161 >= `INH(p158)) ? `INH(p158) : f161;
        f161 = (f161 >= `INH(p169)) ? `INH(p169) : f161;
        f162 = 2047;
        f162 = (f162 >= `INH(p171)) ? `INH(p171) : f162;
        f162 = (f162 >= `INH(p172)) ? `INH(p172) : f162;
        f162 = (f162 > p176) ? p176 : f162;
        f163 = 2047;
        f163 = (f163 > p170) ? p170 : f163;
        f163 = (f163 >= `INH(p176)) ? `INH(p176) : f163;
        f164 = 2047;
        f164 = (f164 > p174) ? p174 : f164;
        f164 = (f164 >= `INH(p176)) ? `INH(p176) : f164;
        f165 = 2047;
        f165 = (f165 >= p171/2) ? p171/2 : f165;
        f165 = (f165 >= `INH(p175)) ? `INH(p175) : f165;
        f166 = 2047;
        f166 = (f166 >= `INH(p175)) ? `INH(p175) : f166;
        f166 = (f166 > p178) ? p178 : f166;
        f167 = 2047;
        f167 = (f167 > p171) ? p171 : f167;
        f167 = (f167 >= `INH(p178)) ? `INH(p178) : f167;
        f167 = (f167 > p180) ? p180 : f167;
        f168 = 2047;
        f168 = (f168 >= `INH(p178)) ? `INH(p178) : f168;
        f168 = (f168 > p181) ? p181 : f168;
        f169 = 2047;
        f169 = (f169 > p170) ? p170 : f169;
        f169 = (f169 >= `INH(p180)) ? `INH(p180) : f169;
        f169 = (f169 >= `INH(p181)) ? `INH(p181) : f169;
        f170 = 2047;
        f170 = (f170 > p170) ? p170 : f170;
        f170 = (f170 >= `INH(p179)) ? `INH(p179) : f170;
        f170 = (f170 >= `INH(p181)) ? `INH(p181) : f170;
        f171 = 2047;
        f171 = (f171 >= `INH(p181)) ? `INH(p181) : f171;
        f171 = (f171 > p183) ? p183 : f171;
        f172 = 2047;
        f172 = (f172 > p177) ? p177 : f172;
        f172 = (f172 >= `INH(p183)) ? `INH(p183) : f172;
        f173 = 2047;
        f173 = (f173 >= `INH(p183)) ? `INH(p183) : f173;
        f173 = (f173 > p184) ? p184 : f173;
        f174 = 2047;
        f174 = (f174 > p182) ? p182 : f174;
        f174 = (f174 >= `INH(p184)) ? `INH(p184) : f174;
        f175 = 2047;
        f175 = (f175 > p172) ? p172 : f175;
        f175 = (f175 > p179) ? p179 : f175;
        f175 = (f175 >= `INH(p180)) ? `INH(p180) : f175;
        f175 = (f175 >= `INH(p184)) ? `INH(p184) : f175;
        f176 = 2047;
        f176 = (f176 > p172) ? p172 : f176;
        f176 = (f176 >= `INH(p179)) ? `INH(p179) : f176;
        f176 = (f176 >= `INH(p184)) ? `INH(p184) : f176;
        f177 = 2047;
        f177 = (f177 > p28) ? p28 : f177;
        f177 = (f177 >= `INH(p186)) ? `INH(p186) : f177;
        f178 = 2047;
        f178 = (f178 > p185) ? p185 : f178;
        f178 = (f178 >= `INH(p187)) ? `INH(p187) : f178;
        f179 = 2047;
        f179 = (f179 >= `INH(p28)) ? `INH(p28) : f179;
        f179 = (f179 >= `INH(p186)) ? `INH(p186) : f179;
        f179 = (f179 > p187) ? p187 : f179;
        f180 = 2047;
        f180 = (f180 >= `INH(p185)) ? `INH(p185) : f180;
        f180 = (f180 >= `INH(p187)) ? `INH(p187) : f180;
        f180 = (f180 > p188) ? p188 : f180;
        f181 = 2047;
        f181 = (f181 > p29) ? p29 : f181;
        f181 = (f181 >= `INH(p190)) ? `INH(p190) : f181;
        f182 = 2047;
        f182 = (f182 > p189) ? p189 : f182;
        f182 = (f182 >= `INH(p191)) ? `INH(p191) : f182;
        f183 = 2047;
        f183 = (f183 >= `INH(p29)) ? `INH(p29) : f183;
        f183 = (f183 >= `INH(p190)) ? `INH(p190) : f183;
        f183 = (f183 > p191) ? p191 : f183;
        f184 = 2047;
        f184 = (f184 >= `INH(p189)) ? `INH(p189) : f184;
        f184 = (f184 >= `INH(p191)) ? `INH(p191) : f184;
        f184 = (f184 > p192) ? p192 : f184;
        f185 = 2047;
        f185 = (f185 >= `INH(p24)) ? `INH(p24) : f185;
        f185 = (f185 > p186) ? p186 : f185;
        f185 = (f185 > p190) ? p190 : f185;
        f186 = 2047;
        f186 = (f186 > p172) ? p172 : f186;
        f186 = (f186 >= `INH(p188)) ? `INH(p188) : f186;
        f186 = (f186 >= `INH(p192)) ? `INH(p192) : f186;
        f187 = 2047;
        f187 = (f187 > p173) ? p173 : f187;
        f187 = (f187 >= `INH(p193)) ? `INH(p193) : f187;
        f188 = 2047;
        f188 = (f188 > p30) ? p30 : f188;
        f188 = (f188 >= `INH(p174)) ? `INH(p174) : f188;
        f189 = 2047;
        f189 = (f189 >= `INH(p30)) ? `INH(p30) : f189;
        f189 = (f189 >= `INH(p174)) ? `INH(p174) : f189;
        f189 = (f189 > p193) ? p193 : f189;
        f190 = 2047;
        f190 = (f190 > p25) ? p25 : f190;
        f190 = (f190 >= `INH(p173)) ? `INH(p173) : f190;
        f190 = (f190 >= `INH(p193)) ? `INH(p193) : f190;
        f191 = 2047;
        f191 = (f191 >= `INH(p195)) ? `INH(p195) : f191;
        f191 = (f191 >= `INH(p196)) ? `INH(p196) : f191;
        f191 = (f191 > p200) ? p200 : f191;
        f192 = 2047;
        f192 = (f192 > p194) ? p194 : f192;
        f192 = (f192 >= `INH(p200)) ? `INH(p200) : f192;
        f193 = 2047;
        f193 = (f193 > p198) ? p198 : f193;
        f193 = (f193 >= `INH(p200)) ? `INH(p200) : f193;
        f194 = 2047;
        f194 = (f194 >= p195/2) ? p195/2 : f194;
        f194 = (f194 >= `INH(p199)) ? `INH(p199) : f194;
        f195 = 2047;
        f195 = (f195 >= `INH(p199)) ? `INH(p199) : f195;
        f195 = (f195 > p202) ? p202 : f195;
        f196 = 2047;
        f196 = (f196 > p195) ? p195 : f196;
        f196 = (f196 >= `INH(p202)) ? `INH(p202) : f196;
        f196 = (f196 > p204) ? p204 : f196;
        f197 = 2047;
        f197 = (f197 >= `INH(p202)) ? `INH(p202) : f197;
        f197 = (f197 > p205) ? p205 : f197;
        f198 = 2047;
        f198 = (f198 > p194) ? p194 : f198;
        f198 = (f198 >= `INH(p204)) ? `INH(p204) : f198;
        f198 = (f198 >= `INH(p205)) ? `INH(p205) : f198;
        f199 = 2047;
        f199 = (f199 > p194) ? p194 : f199;
        f199 = (f199 >= `INH(p203)) ? `INH(p203) : f199;
        f199 = (f199 >= `INH(p205)) ? `INH(p205) : f199;
        f200 = 2047;
        f200 = (f200 >= `INH(p205)) ? `INH(p205) : f200;
        f200 = (f200 > p207) ? p207 : f200;
        f201 = 2047;
        f201 = (f201 > p201) ? p201 : f201;
        f201 = (f201 >= `INH(p207)) ? `INH(p207) : f201;
        f202 = 2047;
        f202 = (f202 >= `INH(p207)) ? `INH(p207) : f202;
        f202 = (f202 > p208) ? p208 : f202;
        f203 = 2047;
        f203 = (f203 > p206) ? p206 : f203;
        f203 = (f203 >= `INH(p208)) ? `INH(p208) : f203;
        f204 = 2047;
        f204 = (f204 > p196) ? p196 : f204;
        f204 = (f204 > p203) ? p203 : f204;
        f204 = (f204 >= `INH(p204)) ? `INH(p204) : f204;
        f204 = (f204 >= `INH(p208)) ? `INH(p208) : f204;
        f205 = 2047;
        f205 = (f205 > p196) ? p196 : f205;
        f205 = (f205 >= `INH(p203)) ? `INH(p203) : f205;
        f205 = (f205 >= `INH(p208)) ? `INH(p208) : f205;
        f206 = 2047;
        f206 = (f206 > p31) ? p31 : f206;
        f206 = (f206 >= `INH(p210)) ? `INH(p210) : f206;
        f207 = 2047;
        f207 = (f207 > p209) ? p209 : f207;
        f207 = (f207 >= `INH(p211)) ? `INH(p211) : f207;
        f208 = 2047;
        f208 = (f208 >= `INH(p31)) ? `INH(p31) : f208;
        f208 = (f208 >= `INH(p210)) ? `INH(p210) : f208;
        f208 = (f208 > p211) ? p211 : f208;
        f209 = 2047;
        f209 = (f209 >= `INH(p209)) ? `INH(p209) : f209;
        f209 = (f209 >= `INH(p211)) ? `INH(p211) : f209;
        f209 = (f209 > p212) ? p212 : f209;
        f210 = 2047;
        f210 = (f210 > p32) ? p32 : f210;
        f210 = (f210 >= `INH(p214)) ? `INH(p214) : f210;
        f211 = 2047;
        f211 = (f211 > p213) ? p213 : f211;
        f211 = (f211 >= `INH(p215)) ? `INH(p215) : f211;
        f212 = 2047;
        f212 = (f212 >= `INH(p32)) ? `INH(p32) : f212;
        f212 = (f212 >= `INH(p214)) ? `INH(p214) : f212;
        f212 = (f212 > p215) ? p215 : f212;
        f213 = 2047;
        f213 = (f213 >= `INH(p213)) ? `INH(p213) : f213;
        f213 = (f213 >= `INH(p215)) ? `INH(p215) : f213;
        f213 = (f213 > p216) ? p216 : f213;
        f214 = 2047;
        f214 = (f214 >= `INH(p25)) ? `INH(p25) : f214;
        f214 = (f214 > p210) ? p210 : f214;
        f214 = (f214 > p214) ? p214 : f214;
        f215 = 2047;
        f215 = (f215 > p196) ? p196 : f215;
        f215 = (f215 >= `INH(p212)) ? `INH(p212) : f215;
        f215 = (f215 >= `INH(p216)) ? `INH(p216) : f215;
        f216 = 2047;
        f216 = (f216 > p197) ? p197 : f216;
        f216 = (f216 >= `INH(p217)) ? `INH(p217) : f216;
        f217 = 2047;
        f217 = (f217 > p33) ? p33 : f217;
        f217 = (f217 >= `INH(p198)) ? `INH(p198) : f217;
        f218 = 2047;
        f218 = (f218 >= `INH(p33)) ? `INH(p33) : f218;
        f218 = (f218 >= `INH(p198)) ? `INH(p198) : f218;
        f218 = (f218 > p217) ? p217 : f218;
        f219 = 2047;
        f219 = (f219 > p26) ? p26 : f219;
        f219 = (f219 >= `INH(p197)) ? `INH(p197) : f219;
        f219 = (f219 >= `INH(p217)) ? `INH(p217) : f219;
        f220 = 2047;
        f220 = (f220 > p219) ? p219 : f220;
        f220 = (f220 >= `INH(p221)) ? `INH(p221) : f220;
        f221 = 2047;
        f221 = (f221 >= `INH(p218)) ? `INH(p218) : f221;
        f221 = (f221 >= `INH(p219)) ? `INH(p219) : f221;
        f221 = (f221 >= `INH(p221)) ? `INH(p221) : f221;
        f221 = (f221 > p222) ? p222 : f221;
        f222 = 2047;
        f222 = (f222 > p30) ? p30 : f222;
        f222 = (f222 >= `INH(p224)) ? `INH(p224) : f222;
        f223 = 2047;
        f223 = (f223 > p223) ? p223 : f223;
        f223 = (f223 >= `INH(p225)) ? `INH(p225) : f223;
        f224 = 2047;
        f224 = (f224 >= `INH(p30)) ? `INH(p30) : f224;
        f224 = (f224 >= `INH(p224)) ? `INH(p224) : f224;
        f224 = (f224 > p225) ? p225 : f224;
        f225 = 2047;
        f225 = (f225 >= `INH(p223)) ? `INH(p223) : f225;
        f225 = (f225 >= `INH(p225)) ? `INH(p225) : f225;
        f225 = (f225 > p226) ? p226 : f225;
        f226 = 2047;
        f226 = (f226 > p33) ? p33 : f226;
        f226 = (f226 >= `INH(p228)) ? `INH(p228) : f226;
        f227 = 2047;
        f227 = (f227 > p227) ? p227 : f227;
        f227 = (f227 >= `INH(p229)) ? `INH(p229) : f227;
        f228 = 2047;
        f228 = (f228 >= `INH(p33)) ? `INH(p33) : f228;
        f228 = (f228 >= `INH(p228)) ? `INH(p228) : f228;
        f228 = (f228 > p229) ? p229 : f228;
        f229 = 2047;
        f229 = (f229 >= `INH(p227)) ? `INH(p227) : f229;
        f229 = (f229 >= `INH(p229)) ? `INH(p229) : f229;
        f229 = (f229 > p230) ? p230 : f229;
        f230 = 2047;
        f230 = (f230 >= `INH(p26)) ? `INH(p26) : f230;
        f230 = (f230 > p224) ? p224 : f230;
        f230 = (f230 > p228) ? p228 : f230;
        f231 = 2047;
        f231 = (f231 > p221) ? p221 : f231;
        f231 = (f231 >= `INH(p226)) ? `INH(p226) : f231;
        f231 = (f231 >= `INH(p230)) ? `INH(p230) : f231;
        f232 = 2047;
        f232 = (f232 > p220) ? p220 : f232;
        f232 = (f232 >= `INH(p231)) ? `INH(p231) : f232;
        f233 = 2047;
        f233 = (f233 > p34) ? p34 : f233;
        f233 = (f233 >= `INH(p222)) ? `INH(p222) : f233;
        f234 = 2047;
        f234 = (f234 >= `INH(p34)) ? `INH(p34) : f234;
        f234 = (f234 >= `INH(p222)) ? `INH(p222) : f234;
        f234 = (f234 > p231) ? p231 : f234;
        f235 = 2047;
        f235 = (f235 > p27) ? p27 : f235;
        f235 = (f235 >= `INH(p220)) ? `INH(p220) : f235;
        f235 = (f235 >= `INH(p231)) ? `INH(p231) : f235;
        f236 = 2047;
        f236 = (f236 >= `INH(p233)) ? `INH(p233) : f236;
        f236 = (f236 >= `INH(p234)) ? `INH(p234) : f236;
        f236 = (f236 > p238) ? p238 : f236;
        f237 = 2047;
        f237 = (f237 > p232) ? p232 : f237;
        f237 = (f237 >= `INH(p238)) ? `INH(p238) : f237;
        f238 = 2047;
        f238 = (f238 > p236) ? p236 : f238;
        f238 = (f238 >= `INH(p238)) ? `INH(p238) : f238;
        f239 = 2047;
        f239 = (f239 >= p233/2) ? p233/2 : f239;
        f239 = (f239 >= `INH(p237)) ? `INH(p237) : f239;
        f240 = 2047;
        f240 = (f240 >= `INH(p237)) ? `INH(p237) : f240;
        f240 = (f240 > p240) ? p240 : f240;
        f241 = 2047;
        f241 = (f241 > p233) ? p233 : f241;
        f241 = (f241 >= `INH(p240)) ? `INH(p240) : f241;
        f241 = (f241 > p242) ? p242 : f241;
        f242 = 2047;
        f242 = (f242 >= `INH(p240)) ? `INH(p240) : f242;
        f242 = (f242 > p243) ? p243 : f242;
        f243 = 2047;
        f243 = (f243 > p232) ? p232 : f243;
        f243 = (f243 >= `INH(p242)) ? `INH(p242) : f243;
        f243 = (f243 >= `INH(p243)) ? `INH(p243) : f243;
        f244 = 2047;
        f244 = (f244 > p232) ? p232 : f244;
        f244 = (f244 >= `INH(p241)) ? `INH(p241) : f244;
        f244 = (f244 >= `INH(p243)) ? `INH(p243) : f244;
        f245 = 2047;
        f245 = (f245 >= `INH(p243)) ? `INH(p243) : f245;
        f245 = (f245 > p245) ? p245 : f245;
        f246 = 2047;
        f246 = (f246 > p239) ? p239 : f246;
        f246 = (f246 >= `INH(p245)) ? `INH(p245) : f246;
        f247 = 2047;
        f247 = (f247 >= `INH(p245)) ? `INH(p245) : f247;
        f247 = (f247 > p246) ? p246 : f247;
        f248 = 2047;
        f248 = (f248 > p244) ? p244 : f248;
        f248 = (f248 >= `INH(p246)) ? `INH(p246) : f248;
        f249 = 2047;
        f249 = (f249 > p234) ? p234 : f249;
        f249 = (f249 > p241) ? p241 : f249;
        f249 = (f249 >= `INH(p242)) ? `INH(p242) : f249;
        f249 = (f249 >= `INH(p246)) ? `INH(p246) : f249;
        f250 = 2047;
        f250 = (f250 > p234) ? p234 : f250;
        f250 = (f250 >= `INH(p241)) ? `INH(p241) : f250;
        f250 = (f250 >= `INH(p246)) ? `INH(p246) : f250;
        f251 = 2047;
        f251 = (f251 > p39) ? p39 : f251;
        f251 = (f251 >= `INH(p248)) ? `INH(p248) : f251;
        f252 = 2047;
        f252 = (f252 > p247) ? p247 : f252;
        f252 = (f252 >= `INH(p249)) ? `INH(p249) : f252;
        f253 = 2047;
        f253 = (f253 >= `INH(p39)) ? `INH(p39) : f253;
        f253 = (f253 >= `INH(p248)) ? `INH(p248) : f253;
        f253 = (f253 > p249) ? p249 : f253;
        f254 = 2047;
        f254 = (f254 >= `INH(p247)) ? `INH(p247) : f254;
        f254 = (f254 >= `INH(p249)) ? `INH(p249) : f254;
        f254 = (f254 > p250) ? p250 : f254;
        f255 = 2047;
        f255 = (f255 > p40) ? p40 : f255;
        f255 = (f255 >= `INH(p252)) ? `INH(p252) : f255;
        f256 = 2047;
        f256 = (f256 > p251) ? p251 : f256;
        f256 = (f256 >= `INH(p253)) ? `INH(p253) : f256;
        f257 = 2047;
        f257 = (f257 >= `INH(p40)) ? `INH(p40) : f257;
        f257 = (f257 >= `INH(p252)) ? `INH(p252) : f257;
        f257 = (f257 > p253) ? p253 : f257;
        f258 = 2047;
        f258 = (f258 >= `INH(p251)) ? `INH(p251) : f258;
        f258 = (f258 >= `INH(p253)) ? `INH(p253) : f258;
        f258 = (f258 > p254) ? p254 : f258;
        f259 = 2047;
        f259 = (f259 >= `INH(p35)) ? `INH(p35) : f259;
        f259 = (f259 > p248) ? p248 : f259;
        f259 = (f259 > p252) ? p252 : f259;
        f260 = 2047;
        f260 = (f260 > p234) ? p234 : f260;
        f260 = (f260 >= `INH(p250)) ? `INH(p250) : f260;
        f260 = (f260 >= `INH(p254)) ? `INH(p254) : f260;
        f261 = 2047;
        f261 = (f261 > p235) ? p235 : f261;
        f261 = (f261 >= `INH(p255)) ? `INH(p255) : f261;
        f262 = 2047;
        f262 = (f262 > p41) ? p41 : f262;
        f262 = (f262 >= `INH(p236)) ? `INH(p236) : f262;
        f263 = 2047;
        f263 = (f263 >= `INH(p41)) ? `INH(p41) : f263;
        f263 = (f263 >= `INH(p236)) ? `INH(p236) : f263;
        f263 = (f263 > p255) ? p255 : f263;
        f264 = 2047;
        f264 = (f264 > p36) ? p36 : f264;
        f264 = (f264 >= `INH(p235)) ? `INH(p235) : f264;
        f264 = (f264 >= `INH(p255)) ? `INH(p255) : f264;
        f265 = 2047;
        f265 = (f265 >= `INH(p257)) ? `INH(p257) : f265;
        f265 = (f265 >= `INH(p258)) ? `INH(p258) : f265;
        f265 = (f265 > p262) ? p262 : f265;
        f266 = 2047;
        f266 = (f266 > p256) ? p256 : f266;
        f266 = (f266 >= `INH(p262)) ? `INH(p262) : f266;
        f267 = 2047;
        f267 = (f267 > p260) ? p260 : f267;
        f267 = (f267 >= `INH(p262)) ? `INH(p262) : f267;
        f268 = 2047;
        f268 = (f268 >= p257/2) ? p257/2 : f268;
        f268 = (f268 >= `INH(p261)) ? `INH(p261) : f268;
        f269 = 2047;
        f269 = (f269 >= `INH(p261)) ? `INH(p261) : f269;
        f269 = (f269 > p264) ? p264 : f269;
        f270 = 2047;
        f270 = (f270 > p257) ? p257 : f270;
        f270 = (f270 >= `INH(p264)) ? `INH(p264) : f270;
        f270 = (f270 > p266) ? p266 : f270;
        f271 = 2047;
        f271 = (f271 >= `INH(p264)) ? `INH(p264) : f271;
        f271 = (f271 > p267) ? p267 : f271;
        f272 = 2047;
        f272 = (f272 > p256) ? p256 : f272;
        f272 = (f272 >= `INH(p266)) ? `INH(p266) : f272;
        f272 = (f272 >= `INH(p267)) ? `INH(p267) : f272;
        f273 = 2047;
        f273 = (f273 > p256) ? p256 : f273;
        f273 = (f273 >= `INH(p265)) ? `INH(p265) : f273;
        f273 = (f273 >= `INH(p267)) ? `INH(p267) : f273;
        f274 = 2047;
        f274 = (f274 >= `INH(p267)) ? `INH(p267) : f274;
        f274 = (f274 > p269) ? p269 : f274;
        f275 = 2047;
        f275 = (f275 > p263) ? p263 : f275;
        f275 = (f275 >= `INH(p269)) ? `INH(p269) : f275;
        f276 = 2047;
        f276 = (f276 >= `INH(p269)) ? `INH(p269) : f276;
        f276 = (f276 > p270) ? p270 : f276;
        f277 = 2047;
        f277 = (f277 > p268) ? p268 : f277;
        f277 = (f277 >= `INH(p270)) ? `INH(p270) : f277;
        f278 = 2047;
        f278 = (f278 > p258) ? p258 : f278;
        f278 = (f278 > p265) ? p265 : f278;
        f278 = (f278 >= `INH(p266)) ? `INH(p266) : f278;
        f278 = (f278 >= `INH(p270)) ? `INH(p270) : f278;
        f279 = 2047;
        f279 = (f279 > p258) ? p258 : f279;
        f279 = (f279 >= `INH(p265)) ? `INH(p265) : f279;
        f279 = (f279 >= `INH(p270)) ? `INH(p270) : f279;
        f280 = 2047;
        f280 = (f280 > p42) ? p42 : f280;
        f280 = (f280 >= `INH(p272)) ? `INH(p272) : f280;
        f281 = 2047;
        f281 = (f281 > p271) ? p271 : f281;
        f281 = (f281 >= `INH(p273)) ? `INH(p273) : f281;
        f282 = 2047;
        f282 = (f282 >= `INH(p42)) ? `INH(p42) : f282;
        f282 = (f282 >= `INH(p272)) ? `INH(p272) : f282;
        f282 = (f282 > p273) ? p273 : f282;
        f283 = 2047;
        f283 = (f283 >= `INH(p271)) ? `INH(p271) : f283;
        f283 = (f283 >= `INH(p273)) ? `INH(p273) : f283;
        f283 = (f283 > p274) ? p274 : f283;
        f284 = 2047;
        f284 = (f284 > p43) ? p43 : f284;
        f284 = (f284 >= `INH(p276)) ? `INH(p276) : f284;
        f285 = 2047;
        f285 = (f285 > p275) ? p275 : f285;
        f285 = (f285 >= `INH(p277)) ? `INH(p277) : f285;
        f286 = 2047;
        f286 = (f286 >= `INH(p43)) ? `INH(p43) : f286;
        f286 = (f286 >= `INH(p276)) ? `INH(p276) : f286;
        f286 = (f286 > p277) ? p277 : f286;
        f287 = 2047;
        f287 = (f287 >= `INH(p275)) ? `INH(p275) : f287;
        f287 = (f287 >= `INH(p277)) ? `INH(p277) : f287;
        f287 = (f287 > p278) ? p278 : f287;
        f288 = 2047;
        f288 = (f288 >= `INH(p36)) ? `INH(p36) : f288;
        f288 = (f288 > p272) ? p272 : f288;
        f288 = (f288 > p276) ? p276 : f288;
        f289 = 2047;
        f289 = (f289 > p258) ? p258 : f289;
        f289 = (f289 >= `INH(p274)) ? `INH(p274) : f289;
        f289 = (f289 >= `INH(p278)) ? `INH(p278) : f289;
        f290 = 2047;
        f290 = (f290 > p259) ? p259 : f290;
        f290 = (f290 >= `INH(p279)) ? `INH(p279) : f290;
        f291 = 2047;
        f291 = (f291 > p44) ? p44 : f291;
        f291 = (f291 >= `INH(p260)) ? `INH(p260) : f291;
        f292 = 2047;
        f292 = (f292 >= `INH(p44)) ? `INH(p44) : f292;
        f292 = (f292 >= `INH(p260)) ? `INH(p260) : f292;
        f292 = (f292 > p279) ? p279 : f292;
        f293 = 2047;
        f293 = (f293 > p37) ? p37 : f293;
        f293 = (f293 >= `INH(p259)) ? `INH(p259) : f293;
        f293 = (f293 >= `INH(p279)) ? `INH(p279) : f293;
        f294 = 2047;
        f294 = (f294 > p281) ? p281 : f294;
        f294 = (f294 >= `INH(p283)) ? `INH(p283) : f294;
        f295 = 2047;
        f295 = (f295 >= `INH(p280)) ? `INH(p280) : f295;
        f295 = (f295 >= `INH(p281)) ? `INH(p281) : f295;
        f295 = (f295 >= `INH(p283)) ? `INH(p283) : f295;
        f295 = (f295 > p284) ? p284 : f295;
        f296 = 2047;
        f296 = (f296 > p41) ? p41 : f296;
        f296 = (f296 >= `INH(p286)) ? `INH(p286) : f296;
        f297 = 2047;
        f297 = (f297 > p285) ? p285 : f297;
        f297 = (f297 >= `INH(p287)) ? `INH(p287) : f297;
        f298 = 2047;
        f298 = (f298 >= `INH(p41)) ? `INH(p41) : f298;
        f298 = (f298 >= `INH(p286)) ? `INH(p286) : f298;
        f298 = (f298 > p287) ? p287 : f298;
        f299 = 2047;
        f299 = (f299 >= `INH(p285)) ? `INH(p285) : f299;
        f299 = (f299 >= `INH(p287)) ? `INH(p287) : f299;
        f299 = (f299 > p288) ? p288 : f299;
        f300 = 2047;
        f300 = (f300 > p44) ? p44 : f300;
        f300 = (f300 >= `INH(p290)) ? `INH(p290) : f300;
        f301 = 2047;
        f301 = (f301 > p289) ? p289 : f301;
        f301 = (f301 >= `INH(p291)) ? `INH(p291) : f301;
        f302 = 2047;
        f302 = (f302 >= `INH(p44)) ? `INH(p44) : f302;
        f302 = (f302 >= `INH(p290)) ? `INH(p290) : f302;
        f302 = (f302 > p291) ? p291 : f302;
        f303 = 2047;
        f303 = (f303 >= `INH(p289)) ? `INH(p289) : f303;
        f303 = (f303 >= `INH(p291)) ? `INH(p291) : f303;
        f303 = (f303 > p292) ? p292 : f303;
        f304 = 2047;
        f304 = (f304 >= `INH(p37)) ? `INH(p37) : f304;
        f304 = (f304 > p286) ? p286 : f304;
        f304 = (f304 > p290) ? p290 : f304;
        f305 = 2047;
        f305 = (f305 > p283) ? p283 : f305;
        f305 = (f305 >= `INH(p288)) ? `INH(p288) : f305;
        f305 = (f305 >= `INH(p292)) ? `INH(p292) : f305;
        f306 = 2047;
        f306 = (f306 > p282) ? p282 : f306;
        f306 = (f306 >= `INH(p293)) ? `INH(p293) : f306;
        f307 = 2047;
        f307 = (f307 > p45) ? p45 : f307;
        f307 = (f307 >= `INH(p284)) ? `INH(p284) : f307;
        f308 = 2047;
        f308 = (f308 >= `INH(p45)) ? `INH(p45) : f308;
        f308 = (f308 >= `INH(p284)) ? `INH(p284) : f308;
        f308 = (f308 > p293) ? p293 : f308;
        f309 = 2047;
        f309 = (f309 > p38) ? p38 : f309;
        f309 = (f309 >= `INH(p282)) ? `INH(p282) : f309;
        f309 = (f309 >= `INH(p293)) ? `INH(p293) : f309;
        if(f14>0)
                f2 = 0;
        if(f15>0)
                f16 = 0;
        if(f17>0)
                f18 = 0;
        if(f19>0)
                f20 = 0;
        if(f21>0)
                f23 = 0;
        if(f22>0)
                f23 = 0;
        if(f24>0)
                f25 = 0;
        if(f26>0)
                f27 = 0;
        if(f26>0)
                f28 = 0;
        if(f43>0)
                f3 = 0;
        if(f44>0)
                f45 = 0;
        if(f46>0)
                f47 = 0;
        if(f48>0)
                f49 = 0;
        if(f50>0)
                f52 = 0;
        if(f51>0)
                f52 = 0;
        if(f53>0)
                f54 = 0;
        if(f55>0)
                f56 = 0;
        if(f55>0)
                f57 = 0;
        if(f88>0)
                f5 = 0;
        if(f89>0)
                f90 = 0;
        if(f91>0)
                f92 = 0;
        if(f93>0)
                f94 = 0;
        if(f95>0)
                f97 = 0;
        if(f96>0)
                f97 = 0;
        if(f98>0)
                f99 = 0;
        if(f100>0)
                f101 = 0;
        if(f100>0)
                f102 = 0;
        if(f117>0)
                f6 = 0;
        if(f118>0)
                f119 = 0;
        if(f120>0)
                f121 = 0;
        if(f122>0)
                f123 = 0;
        if(f124>0)
                f126 = 0;
        if(f125>0)
                f126 = 0;
        if(f127>0)
                f128 = 0;
        if(f129>0)
                f130 = 0;
        if(f129>0)
                f131 = 0;
        if(f162>0)
                f8 = 0;
        if(f163>0)
                f164 = 0;
        if(f165>0)
                f166 = 0;
        if(f167>0)
                f168 = 0;
        if(f169>0)
                f171 = 0;
        if(f170>0)
                f171 = 0;
        if(f172>0)
                f173 = 0;
        if(f174>0)
                f175 = 0;
        if(f174>0)
                f176 = 0;
        if(f191>0)
                f9 = 0;
        if(f192>0)
                f193 = 0;
        if(f194>0)
                f195 = 0;
        if(f196>0)
                f197 = 0;
        if(f198>0)
                f200 = 0;
        if(f199>0)
                f200 = 0;
        if(f201>0)
                f202 = 0;
        if(f203>0)
                f204 = 0;
        if(f203>0)
                f205 = 0;
        if(f236>0)
                f11 = 0;
        if(f237>0)
                f238 = 0;
        if(f239>0)
                f240 = 0;
        if(f241>0)
                f242 = 0;
        if(f243>0)
                f245 = 0;
        if(f244>0)
                f245 = 0;
        if(f246>0)
                f247 = 0;
        if(f248>0)
                f249 = 0;
        if(f248>0)
                f250 = 0;
        if(f265>0)
                f12 = 0;
        if(f266>0)
                f267 = 0;
        if(f268>0)
                f269 = 0;
        if(f270>0)
                f271 = 0;
        if(f272>0)
                f274 = 0;
        if(f273>0)
                f274 = 0;
        if(f275>0)
                f276 = 0;
        if(f277>0)
                f278 = 0;
        if(f277>0)
                f279 = 0;
        tf = (f0>0)?1:(f1>0)?2:(f2>0)?3:(f3>0)?4:(f4>0)?5:(f5>0)?6:(f6>0)?7:(f7>0)?8:(f8>0)?9:(f9>0)?10:(f10>0)?11:(f11>0)?12:(f12>0)?13:(f13>0)?14:(f14>0)?15:(f15>0)?16:(f16>0)?17:(f17>0)?18:(f18>0)?19:(f19>0)?20:(f20>0)?21:(f21>0)?22:(f22>0)?23:(f23>0)?24:(f24>0)?25:(f25>0)?26:(f26>0)?27:(f27>0)?28:(f28>0)?29:(f29>0)?30:(f30>0)?31:(f31>0)?32:(f32>0)?33:(f33>0)?34:(f34>0)?35:(f35>0)?36:(f36>0)?37:(f37>0)?38:(f38>0)?39:(f39>0)?40:(f40>0)?41:(f41>0)?42:(f42>0)?43:(f43>0)?44:(f44>0)?45:(f45>0)?46:(f46>0)?47:(f47>0)?48:(f48>0)?49:(f49>0)?50:(f50>0)?51:(f51>0)?52:(f52>0)?53:(f53>0)?54:(f54>0)?55:(f55>0)?56:(f56>0)?57:(f57>0)?58:(f58>0)?59:(f59>0)?60:(f60>0)?61:(f61>0)?62:(f62>0)?63:(f63>0)?64:(f64>0)?65:(f65>0)?66:(f66>0)?67:(f67>0)?68:(f68>0)?69:(f69>0)?70:(f70>0)?71:(f71>0)?72:(f72>0)?73:(f73>0)?74:(f74>0)?75:(f75>0)?76:(f76>0)?77:(f77>0)?78:(f78>0)?79:(f79>0)?80:(f80>0)?81:(f81>0)?82:(f82>0)?83:(f83>0)?84:(f84>0)?85:(f85>0)?86:(f86>0)?87:(f87>0)?88:(f88>0)?89:(f89>0)?90:(f90>0)?91:(f91>0)?92:(f92>0)?93:(f93>0)?94:(f94>0)?95:(f95>0)?96:(f96>0)?97:(f97>0)?98:(f98>0)?99:(f99>0)?100:(f100>0)?101:(f101>0)?102:(f102>0)?103:(f103>0)?104:(f104>0)?105:(f105>0)?106:(f106>0)?107:(f107>0)?108:(f108>0)?109:(f109>0)?110:(f110>0)?111:(f111>0)?112:(f112>0)?113:(f113>0)?114:(f114>0)?115:(f115>0)?116:(f116>0)?117:(f117>0)?118:(f118>0)?119:(f119>0)?120:(f120>0)?121:(f121>0)?122:(f122>0)?123:(f123>0)?124:(f124>0)?125:(f125>0)?126:(f126>0)?127:(f127>0)?128:(f128>0)?129:(f129>0)?130:(f130>0)?131:(f131>0)?132:(f132>0)?133:(f133>0)?134:(f134>0)?135:(f135>0)?136:(f136>0)?137:(f137>0)?138:(f138>0)?139:(f139>0)?140:(f140>0)?141:(f141>0)?142:(f142>0)?143:(f143>0)?144:(f144>0)?145:(f145>0)?146:(f146>0)?147:(f147>0)?148:(f148>0)?149:(f149>0)?150:(f150>0)?151:(f151>0)?152:(f152>0)?153:(f153>0)?154:(f154>0)?155:(f155>0)?156:(f156>0)?157:(f157>0)?158:(f158>0)?159:(f159>0)?160:(f160>0)?161:(f161>0)?162:(f162>0)?163:(f163>0)?164:(f164>0)?165:(f165>0)?166:(f166>0)?167:(f167>0)?168:(f168>0)?169:(f169>0)?170:(f170>0)?171:(f171>0)?172:(f172>0)?173:(f173>0)?174:(f174>0)?175:(f175>0)?176:(f176>0)?177:(f177>0)?178:(f178>0)?179:(f179>0)?180:(f180>0)?181:(f181>0)?182:(f182>0)?183:(f183>0)?184:(f184>0)?185:(f185>0)?186:(f186>0)?187:(f187>0)?188:(f188>0)?189:(f189>0)?190:(f190>0)?191:(f191>0)?192:(f192>0)?193:(f193>0)?194:(f194>0)?195:(f195>0)?196:(f196>0)?197:(f197>0)?198:(f198>0)?199:(f199>0)?200:(f200>0)?201:(f201>0)?202:(f202>0)?203:(f203>0)?204:(f204>0)?205:(f205>0)?206:(f206>0)?207:(f207>0)?208:(f208>0)?209:(f209>0)?210:(f210>0)?211:(f211>0)?212:(f212>0)?213:(f213>0)?214:(f214>0)?215:(f215>0)?216:(f216>0)?217:(f217>0)?218:(f218>0)?219:(f219>0)?220:(f220>0)?221:(f221>0)?222:(f222>0)?223:(f223>0)?224:(f224>0)?225:(f225>0)?226:(f226>0)?227:(f227>0)?228:(f228>0)?229:(f229>0)?230:(f230>0)?231:(f231>0)?232:(f232>0)?233:(f233>0)?234:(f234>0)?235:(f235>0)?236:(f236>0)?237:(f237>0)?238:(f238>0)?239:(f239>0)?240:(f240>0)?241:(f241>0)?242:(f242>0)?243:(f243>0)?244:(f244>0)?245:(f245>0)?246:(f246>0)?247:(f247>0)?248:(f248>0)?249:(f249>0)?250:(f250>0)?251:(f251>0)?252:(f252>0)?253:(f253>0)?254:(f254>0)?255:(f255>0)?256:(f256>0)?257:(f257>0)?258:(f258>0)?259:(f259>0)?260:(f260>0)?261:(f261>0)?262:(f262>0)?263:(f263>0)?264:(f264>0)?265:(f265>0)?266:(f266>0)?267:(f267>0)?268:(f268>0)?269:(f269>0)?270:(f270>0)?271:(f271>0)?272:(f272>0)?273:(f273>0)?274:(f274>0)?275:(f275>0)?276:(f276>0)?277:(f277>0)?278:(f278>0)?279:(f279>0)?280:(f280>0)?281:(f281>0)?282:(f282>0)?283:(f283>0)?284:(f284>0)?285:(f285>0)?286:(f286>0)?287:(f287>0)?288:(f288>0)?289:(f289>0)?290:(f290>0)?291:(f291>0)?292:(f292>0)?293:(f293>0)?294:(f294>0)?295:(f295>0)?296:(f296>0)?297:(f297>0)?298:(f298>0)?299:(f299>0)?300:(f300>0)?301:(f301>0)?302:(f302>0)?303:(f303>0)?304:(f304>0)?305:(f305>0)?306:(f306>0)?307:(f307>0)?308:(f308>0)?309:(f309>0)?310:0;
        case(tf)
                1: begin
                        tc = f0;
                        p2 = p2 - tc;
                        p13 = p13 - tc;
                        p24 = p24 - tc;
                        p35 = p35 - tc;
                        p0 = p0 + tc;
                end
                2: begin
                        tc = f1;
                        p1 = p1 - tc;
                        p5 = p5 + tc;
                        p16 = p16 + tc;
                        p27 = p27 + tc;
                        p38 = p38 + tc;
                end
                3: begin
                        tc = f2;
                        p51 = p51 - tc;
                        p48 = p48 + tc;
                end
                4: begin
                        tc = f3;
                        p75 = p75 - tc;
                        p72 = p72 + tc;
                end
                5: begin
                        tc = f4;
                        p94 = p94 - tc;
                        p96 = p96 + tc;
                end
                6: begin
                        tc = f5;
                        p113 = p113 - tc;
                        p110 = p110 + tc;
                end
                7: begin
                        tc = f6;
                        p137 = p137 - tc;
                        p134 = p134 + tc;
                end
                8: begin
                        tc = f7;
                        p156 = p156 - tc;
                        p158 = p158 + tc;
                end
                9: begin
                        tc = f8;
                        p175 = p175 - tc;
                        p172 = p172 + tc;
                end
                10: begin
                        tc = f9;
                        p199 = p199 - tc;
                        p196 = p196 + tc;
                end
                11: begin
                        tc = f10;
                        p218 = p218 - tc;
                        p220 = p220 + tc;
                end
                12: begin
                        tc = f11;
                        p237 = p237 - tc;
                        p234 = p234 + tc;
                end
                13: begin
                        tc = f12;
                        p261 = p261 - tc;
                        p258 = p258 + tc;
                end
                14: begin
                        tc = f13;
                        p280 = p280 - tc;
                        p282 = p282 + tc;
                end
                15: begin
                        tc = f14;
                        p52 = p52 - tc;
                        p48 = p48 + tc;
                end
                16: begin
                        tc = f15;
                        p46 = p46 - tc;
                end
                17: begin
                        tc = f16;
                        p50 = p50 - tc;
                        p52 = p52 + tc;
                end
                18: begin
                        tc = f17;
                        p47 = p47 - tc*2;
                        p53 = p53 + tc;
                end
                19: begin
                        tc = f18;
                        p54 = p54 - tc;
                        p51 = p51 + tc;
                end
                20: begin
                        tc = f19;
                        p47 = p47 - tc;
                        p56 = p56 - tc;
                        p55 = p55 + tc;
                end
                21: begin
                        tc = f20;
                        p57 = p57 - tc;
                        p54 = p54 + tc;
                end
                22: begin
                        tc = f21;
                        p46 = p46 - tc;
                        p49 = p49 + tc;
                        p58 = p58 + tc;
                end
                23: begin
                        tc = f22;
                        p46 = p46 - tc;
                        p58 = p58 + tc;
                end
                24: begin
                        tc = f23;
                        p59 = p59 - tc;
                        p57 = p57 + tc;
                end
                25: begin
                        tc = f24;
                        p53 = p53 - tc;
                        p47 = p47 + tc;
                end
                26: begin
                        tc = f25;
                        p60 = p60 - tc;
                        p59 = p59 + tc;
                end
                27: begin
                        tc = f26;
                        p58 = p58 - tc;
                        p46 = p46 + tc*2;
                end
                28: begin
                        tc = f27;
                        p48 = p48 - tc;
                        p55 = p55 - tc;
                        p56 = p56 + tc;
                        p60 = p60 + tc;
                end
                29: begin
                        tc = f28;
                        p48 = p48 - tc;
                        p60 = p60 + tc;
                end
                30: begin
                        tc = f29;
                        p6 = p6 - tc;
                        p46 = p46 + tc;
                        p61 = p61 + tc;
                end
                31: begin
                        tc = f30;
                        p61 = p61 - tc;
                        p6 = p6 + tc;
                end
                32: begin
                        tc = f31;
                        p63 = p63 - tc;
                        p62 = p62 + tc;
                end
                33: begin
                        tc = f32;
                        p64 = p64 - tc;
                        p63 = p63 + tc;
                end
                34: begin
                        tc = f33;
                        p7 = p7 - tc;
                        p47 = p47 + tc;
                        p65 = p65 + tc;
                end
                35: begin
                        tc = f34;
                        p65 = p65 - tc;
                        p7 = p7 + tc;
                end
                36: begin
                        tc = f35;
                        p67 = p67 - tc;
                        p66 = p66 + tc;
                end
                37: begin
                        tc = f36;
                        p68 = p68 - tc;
                        p67 = p67 + tc;
                end
                38: begin
                        tc = f37;
                        p62 = p62 - tc;
                        p66 = p66 - tc;
                        p2 = p2 + tc;
                end
                39: begin
                        tc = f38;
                        p48 = p48 - tc;
                        p64 = p64 + tc;
                        p68 = p68 + tc;
                end
                40: begin
                        tc = f39;
                        p49 = p49 - tc;
                        p8 = p8 + tc;
                end
                41: begin
                        tc = f40;
                        p8 = p8 - tc;
                end
                42: begin
                        tc = f41;
                        p69 = p69 - tc;
                        p50 = p50 + tc;
                end
                43: begin
                        tc = f42;
                        p3 = p3 - tc;
                        p69 = p69 + tc;
                end
                44: begin
                        tc = f43;
                        p76 = p76 - tc;
                        p72 = p72 + tc;
                end
                45: begin
                        tc = f44;
                        p70 = p70 - tc;
                end
                46: begin
                        tc = f45;
                        p74 = p74 - tc;
                        p76 = p76 + tc;
                end
                47: begin
                        tc = f46;
                        p71 = p71 - tc*2;
                        p77 = p77 + tc;
                end
                48: begin
                        tc = f47;
                        p78 = p78 - tc;
                        p75 = p75 + tc;
                end
                49: begin
                        tc = f48;
                        p71 = p71 - tc;
                        p80 = p80 - tc;
                        p79 = p79 + tc;
                end
                50: begin
                        tc = f49;
                        p81 = p81 - tc;
                        p78 = p78 + tc;
                end
                51: begin
                        tc = f50;
                        p70 = p70 - tc;
                        p73 = p73 + tc;
                        p82 = p82 + tc;
                end
                52: begin
                        tc = f51;
                        p70 = p70 - tc;
                        p82 = p82 + tc;
                end
                53: begin
                        tc = f52;
                        p83 = p83 - tc;
                        p81 = p81 + tc;
                end
                54: begin
                        tc = f53;
                        p77 = p77 - tc;
                        p71 = p71 + tc;
                end
                55: begin
                        tc = f54;
                        p84 = p84 - tc;
                        p83 = p83 + tc;
                end
                56: begin
                        tc = f55;
                        p82 = p82 - tc;
                        p70 = p70 + tc*2;
                end
                57: begin
                        tc = f56;
                        p72 = p72 - tc;
                        p79 = p79 - tc;
                        p80 = p80 + tc;
                        p84 = p84 + tc;
                end
                58: begin
                        tc = f57;
                        p72 = p72 - tc;
                        p84 = p84 + tc;
                end
                59: begin
                        tc = f58;
                        p9 = p9 - tc;
                        p70 = p70 + tc;
                        p85 = p85 + tc;
                end
                60: begin
                        tc = f59;
                        p85 = p85 - tc;
                        p9 = p9 + tc;
                end
                61: begin
                        tc = f60;
                        p87 = p87 - tc;
                        p86 = p86 + tc;
                end
                62: begin
                        tc = f61;
                        p88 = p88 - tc;
                        p87 = p87 + tc;
                end
                63: begin
                        tc = f62;
                        p10 = p10 - tc;
                        p71 = p71 + tc;
                        p89 = p89 + tc;
                end
                64: begin
                        tc = f63;
                        p89 = p89 - tc;
                        p10 = p10 + tc;
                end
                65: begin
                        tc = f64;
                        p91 = p91 - tc;
                        p90 = p90 + tc;
                end
                66: begin
                        tc = f65;
                        p92 = p92 - tc;
                        p91 = p91 + tc;
                end
                67: begin
                        tc = f66;
                        p86 = p86 - tc;
                        p90 = p90 - tc;
                        p3 = p3 + tc;
                end
                68: begin
                        tc = f67;
                        p72 = p72 - tc;
                        p88 = p88 + tc;
                        p92 = p92 + tc;
                end
                69: begin
                        tc = f68;
                        p73 = p73 - tc;
                        p11 = p11 + tc;
                end
                70: begin
                        tc = f69;
                        p11 = p11 - tc;
                end
                71: begin
                        tc = f70;
                        p93 = p93 - tc;
                        p74 = p74 + tc;
                end
                72: begin
                        tc = f71;
                        p4 = p4 - tc;
                        p93 = p93 + tc;
                end
                73: begin
                        tc = f72;
                        p95 = p95 - tc;
                        p96 = p96 + tc;
                end
                74: begin
                        tc = f73;
                        p98 = p98 - tc;
                        p97 = p97 + tc;
                end
                75: begin
                        tc = f74;
                        p8 = p8 - tc;
                        p94 = p94 + tc;
                        p99 = p99 + tc;
                end
                76: begin
                        tc = f75;
                        p99 = p99 - tc;
                        p8 = p8 + tc;
                end
                77: begin
                        tc = f76;
                        p101 = p101 - tc;
                        p100 = p100 + tc;
                end
                78: begin
                        tc = f77;
                        p102 = p102 - tc;
                        p101 = p101 + tc;
                end
                79: begin
                        tc = f78;
                        p11 = p11 - tc;
                        p95 = p95 + tc;
                        p103 = p103 + tc;
                end
                80: begin
                        tc = f79;
                        p103 = p103 - tc;
                        p11 = p11 + tc;
                end
                81: begin
                        tc = f80;
                        p105 = p105 - tc;
                        p104 = p104 + tc;
                end
                82: begin
                        tc = f81;
                        p106 = p106 - tc;
                        p105 = p105 + tc;
                end
                83: begin
                        tc = f82;
                        p100 = p100 - tc;
                        p104 = p104 - tc;
                        p4 = p4 + tc;
                end
                84: begin
                        tc = f83;
                        p97 = p97 - tc;
                        p102 = p102 + tc;
                        p106 = p106 + tc;
                end
                85: begin
                        tc = f84;
                        p96 = p96 - tc;
                        p12 = p12 + tc;
                end
                86: begin
                        tc = f85;
                        p12 = p12 - tc;
                end
                87: begin
                        tc = f86;
                        p107 = p107 - tc;
                        p98 = p98 + tc;
                end
                88: begin
                        tc = f87;
                        p5 = p5 - tc;
                        p107 = p107 + tc;
                end
                89: begin
                        tc = f88;
                        p114 = p114 - tc;
                        p110 = p110 + tc;
                end
                90: begin
                        tc = f89;
                        p108 = p108 - tc;
                end
                91: begin
                        tc = f90;
                        p112 = p112 - tc;
                        p114 = p114 + tc;
                end
                92: begin
                        tc = f91;
                        p109 = p109 - tc*2;
                        p115 = p115 + tc;
                end
                93: begin
                        tc = f92;
                        p116 = p116 - tc;
                        p113 = p113 + tc;
                end
                94: begin
                        tc = f93;
                        p109 = p109 - tc;
                        p118 = p118 - tc;
                        p117 = p117 + tc;
                end
                95: begin
                        tc = f94;
                        p119 = p119 - tc;
                        p116 = p116 + tc;
                end
                96: begin
                        tc = f95;
                        p108 = p108 - tc;
                        p111 = p111 + tc;
                        p120 = p120 + tc;
                end
                97: begin
                        tc = f96;
                        p108 = p108 - tc;
                        p120 = p120 + tc;
                end
                98: begin
                        tc = f97;
                        p121 = p121 - tc;
                        p119 = p119 + tc;
                end
                99: begin
                        tc = f98;
                        p115 = p115 - tc;
                        p109 = p109 + tc;
                end
                100: begin
                        tc = f99;
                        p122 = p122 - tc;
                        p121 = p121 + tc;
                end
                101: begin
                        tc = f100;
                        p120 = p120 - tc;
                        p108 = p108 + tc*2;
                end
                102: begin
                        tc = f101;
                        p110 = p110 - tc;
                        p117 = p117 - tc;
                        p118 = p118 + tc;
                        p122 = p122 + tc;
                end
                103: begin
                        tc = f102;
                        p110 = p110 - tc;
                        p122 = p122 + tc;
                end
                104: begin
                        tc = f103;
                        p17 = p17 - tc;
                        p108 = p108 + tc;
                        p123 = p123 + tc;
                end
                105: begin
                        tc = f104;
                        p123 = p123 - tc;
                        p17 = p17 + tc;
                end
                106: begin
                        tc = f105;
                        p125 = p125 - tc;
                        p124 = p124 + tc;
                end
                107: begin
                        tc = f106;
                        p126 = p126 - tc;
                        p125 = p125 + tc;
                end
                108: begin
                        tc = f107;
                        p18 = p18 - tc;
                        p109 = p109 + tc;
                        p127 = p127 + tc;
                end
                109: begin
                        tc = f108;
                        p127 = p127 - tc;
                        p18 = p18 + tc;
                end
                110: begin
                        tc = f109;
                        p129 = p129 - tc;
                        p128 = p128 + tc;
                end
                111: begin
                        tc = f110;
                        p130 = p130 - tc;
                        p129 = p129 + tc;
                end
                112: begin
                        tc = f111;
                        p124 = p124 - tc;
                        p128 = p128 - tc;
                        p13 = p13 + tc;
                end
                113: begin
                        tc = f112;
                        p110 = p110 - tc;
                        p126 = p126 + tc;
                        p130 = p130 + tc;
                end
                114: begin
                        tc = f113;
                        p111 = p111 - tc;
                        p19 = p19 + tc;
                end
                115: begin
                        tc = f114;
                        p19 = p19 - tc;
                end
                116: begin
                        tc = f115;
                        p131 = p131 - tc;
                        p112 = p112 + tc;
                end
                117: begin
                        tc = f116;
                        p14 = p14 - tc;
                        p131 = p131 + tc;
                end
                118: begin
                        tc = f117;
                        p138 = p138 - tc;
                        p134 = p134 + tc;
                end
                119: begin
                        tc = f118;
                        p132 = p132 - tc;
                end
                120: begin
                        tc = f119;
                        p136 = p136 - tc;
                        p138 = p138 + tc;
                end
                121: begin
                        tc = f120;
                        p133 = p133 - tc*2;
                        p139 = p139 + tc;
                end
                122: begin
                        tc = f121;
                        p140 = p140 - tc;
                        p137 = p137 + tc;
                end
                123: begin
                        tc = f122;
                        p133 = p133 - tc;
                        p142 = p142 - tc;
                        p141 = p141 + tc;
                end
                124: begin
                        tc = f123;
                        p143 = p143 - tc;
                        p140 = p140 + tc;
                end
                125: begin
                        tc = f124;
                        p132 = p132 - tc;
                        p135 = p135 + tc;
                        p144 = p144 + tc;
                end
                126: begin
                        tc = f125;
                        p132 = p132 - tc;
                        p144 = p144 + tc;
                end
                127: begin
                        tc = f126;
                        p145 = p145 - tc;
                        p143 = p143 + tc;
                end
                128: begin
                        tc = f127;
                        p139 = p139 - tc;
                        p133 = p133 + tc;
                end
                129: begin
                        tc = f128;
                        p146 = p146 - tc;
                        p145 = p145 + tc;
                end
                130: begin
                        tc = f129;
                        p144 = p144 - tc;
                        p132 = p132 + tc*2;
                end
                131: begin
                        tc = f130;
                        p134 = p134 - tc;
                        p141 = p141 - tc;
                        p142 = p142 + tc;
                        p146 = p146 + tc;
                end
                132: begin
                        tc = f131;
                        p134 = p134 - tc;
                        p146 = p146 + tc;
                end
                133: begin
                        tc = f132;
                        p20 = p20 - tc;
                        p132 = p132 + tc;
                        p147 = p147 + tc;
                end
                134: begin
                        tc = f133;
                        p147 = p147 - tc;
                        p20 = p20 + tc;
                end
                135: begin
                        tc = f134;
                        p149 = p149 - tc;
                        p148 = p148 + tc;
                end
                136: begin
                        tc = f135;
                        p150 = p150 - tc;
                        p149 = p149 + tc;
                end
                137: begin
                        tc = f136;
                        p21 = p21 - tc;
                        p133 = p133 + tc;
                        p151 = p151 + tc;
                end
                138: begin
                        tc = f137;
                        p151 = p151 - tc;
                        p21 = p21 + tc;
                end
                139: begin
                        tc = f138;
                        p153 = p153 - tc;
                        p152 = p152 + tc;
                end
                140: begin
                        tc = f139;
                        p154 = p154 - tc;
                        p153 = p153 + tc;
                end
                141: begin
                        tc = f140;
                        p148 = p148 - tc;
                        p152 = p152 - tc;
                        p14 = p14 + tc;
                end
                142: begin
                        tc = f141;
                        p134 = p134 - tc;
                        p150 = p150 + tc;
                        p154 = p154 + tc;
                end
                143: begin
                        tc = f142;
                        p135 = p135 - tc;
                        p22 = p22 + tc;
                end
                144: begin
                        tc = f143;
                        p22 = p22 - tc;
                end
                145: begin
                        tc = f144;
                        p155 = p155 - tc;
                        p136 = p136 + tc;
                end
                146: begin
                        tc = f145;
                        p15 = p15 - tc;
                        p155 = p155 + tc;
                end
                147: begin
                        tc = f146;
                        p157 = p157 - tc;
                        p158 = p158 + tc;
                end
                148: begin
                        tc = f147;
                        p160 = p160 - tc;
                        p159 = p159 + tc;
                end
                149: begin
                        tc = f148;
                        p19 = p19 - tc;
                        p156 = p156 + tc;
                        p161 = p161 + tc;
                end
                150: begin
                        tc = f149;
                        p161 = p161 - tc;
                        p19 = p19 + tc;
                end
                151: begin
                        tc = f150;
                        p163 = p163 - tc;
                        p162 = p162 + tc;
                end
                152: begin
                        tc = f151;
                        p164 = p164 - tc;
                        p163 = p163 + tc;
                end
                153: begin
                        tc = f152;
                        p22 = p22 - tc;
                        p157 = p157 + tc;
                        p165 = p165 + tc;
                end
                154: begin
                        tc = f153;
                        p165 = p165 - tc;
                        p22 = p22 + tc;
                end
                155: begin
                        tc = f154;
                        p167 = p167 - tc;
                        p166 = p166 + tc;
                end
                156: begin
                        tc = f155;
                        p168 = p168 - tc;
                        p167 = p167 + tc;
                end
                157: begin
                        tc = f156;
                        p162 = p162 - tc;
                        p166 = p166 - tc;
                        p15 = p15 + tc;
                end
                158: begin
                        tc = f157;
                        p159 = p159 - tc;
                        p164 = p164 + tc;
                        p168 = p168 + tc;
                end
                159: begin
                        tc = f158;
                        p158 = p158 - tc;
                        p23 = p23 + tc;
                end
                160: begin
                        tc = f159;
                        p23 = p23 - tc;
                end
                161: begin
                        tc = f160;
                        p169 = p169 - tc;
                        p160 = p160 + tc;
                end
                162: begin
                        tc = f161;
                        p16 = p16 - tc;
                        p169 = p169 + tc;
                end
                163: begin
                        tc = f162;
                        p176 = p176 - tc;
                        p172 = p172 + tc;
                end
                164: begin
                        tc = f163;
                        p170 = p170 - tc;
                end
                165: begin
                        tc = f164;
                        p174 = p174 - tc;
                        p176 = p176 + tc;
                end
                166: begin
                        tc = f165;
                        p171 = p171 - tc*2;
                        p177 = p177 + tc;
                end
                167: begin
                        tc = f166;
                        p178 = p178 - tc;
                        p175 = p175 + tc;
                end
                168: begin
                        tc = f167;
                        p171 = p171 - tc;
                        p180 = p180 - tc;
                        p179 = p179 + tc;
                end
                169: begin
                        tc = f168;
                        p181 = p181 - tc;
                        p178 = p178 + tc;
                end
                170: begin
                        tc = f169;
                        p170 = p170 - tc;
                        p173 = p173 + tc;
                        p182 = p182 + tc;
                end
                171: begin
                        tc = f170;
                        p170 = p170 - tc;
                        p182 = p182 + tc;
                end
                172: begin
                        tc = f171;
                        p183 = p183 - tc;
                        p181 = p181 + tc;
                end
                173: begin
                        tc = f172;
                        p177 = p177 - tc;
                        p171 = p171 + tc;
                end
                174: begin
                        tc = f173;
                        p184 = p184 - tc;
                        p183 = p183 + tc;
                end
                175: begin
                        tc = f174;
                        p182 = p182 - tc;
                        p170 = p170 + tc*2;
                end
                176: begin
                        tc = f175;
                        p172 = p172 - tc;
                        p179 = p179 - tc;
                        p180 = p180 + tc;
                        p184 = p184 + tc;
                end
                177: begin
                        tc = f176;
                        p172 = p172 - tc;
                        p184 = p184 + tc;
                end
                178: begin
                        tc = f177;
                        p28 = p28 - tc;
                        p170 = p170 + tc;
                        p185 = p185 + tc;
                end
                179: begin
                        tc = f178;
                        p185 = p185 - tc;
                        p28 = p28 + tc;
                end
                180: begin
                        tc = f179;
                        p187 = p187 - tc;
                        p186 = p186 + tc;
                end
                181: begin
                        tc = f180;
                        p188 = p188 - tc;
                        p187 = p187 + tc;
                end
                182: begin
                        tc = f181;
                        p29 = p29 - tc;
                        p171 = p171 + tc;
                        p189 = p189 + tc;
                end
                183: begin
                        tc = f182;
                        p189 = p189 - tc;
                        p29 = p29 + tc;
                end
                184: begin
                        tc = f183;
                        p191 = p191 - tc;
                        p190 = p190 + tc;
                end
                185: begin
                        tc = f184;
                        p192 = p192 - tc;
                        p191 = p191 + tc;
                end
                186: begin
                        tc = f185;
                        p186 = p186 - tc;
                        p190 = p190 - tc;
                        p24 = p24 + tc;
                end
                187: begin
                        tc = f186;
                        p172 = p172 - tc;
                        p188 = p188 + tc;
                        p192 = p192 + tc;
                end
                188: begin
                        tc = f187;
                        p173 = p173 - tc;
                        p30 = p30 + tc;
                end
                189: begin
                        tc = f188;
                        p30 = p30 - tc;
                end
                190: begin
                        tc = f189;
                        p193 = p193 - tc;
                        p174 = p174 + tc;
                end
                191: begin
                        tc = f190;
                        p25 = p25 - tc;
                        p193 = p193 + tc;
                end
                192: begin
                        tc = f191;
                        p200 = p200 - tc;
                        p196 = p196 + tc;
                end
                193: begin
                        tc = f192;
                        p194 = p194 - tc;
                end
                194: begin
                        tc = f193;
                        p198 = p198 - tc;
                        p200 = p200 + tc;
                end
                195: begin
                        tc = f194;
                        p195 = p195 - tc*2;
                        p201 = p201 + tc;
                end
                196: begin
                        tc = f195;
                        p202 = p202 - tc;
                        p199 = p199 + tc;
                end
                197: begin
                        tc = f196;
                        p195 = p195 - tc;
                        p204 = p204 - tc;
                        p203 = p203 + tc;
                end
                198: begin
                        tc = f197;
                        p205 = p205 - tc;
                        p202 = p202 + tc;
                end
                199: begin
                        tc = f198;
                        p194 = p194 - tc;
                        p197 = p197 + tc;
                        p206 = p206 + tc;
                end
                200: begin
                        tc = f199;
                        p194 = p194 - tc;
                        p206 = p206 + tc;
                end
                201: begin
                        tc = f200;
                        p207 = p207 - tc;
                        p205 = p205 + tc;
                end
                202: begin
                        tc = f201;
                        p201 = p201 - tc;
                        p195 = p195 + tc;
                end
                203: begin
                        tc = f202;
                        p208 = p208 - tc;
                        p207 = p207 + tc;
                end
                204: begin
                        tc = f203;
                        p206 = p206 - tc;
                        p194 = p194 + tc*2;
                end
                205: begin
                        tc = f204;
                        p196 = p196 - tc;
                        p203 = p203 - tc;
                        p204 = p204 + tc;
                        p208 = p208 + tc;
                end
                206: begin
                        tc = f205;
                        p196 = p196 - tc;
                        p208 = p208 + tc;
                end
                207: begin
                        tc = f206;
                        p31 = p31 - tc;
                        p194 = p194 + tc;
                        p209 = p209 + tc;
                end
                208: begin
                        tc = f207;
                        p209 = p209 - tc;
                        p31 = p31 + tc;
                end
                209: begin
                        tc = f208;
                        p211 = p211 - tc;
                        p210 = p210 + tc;
                end
                210: begin
                        tc = f209;
                        p212 = p212 - tc;
                        p211 = p211 + tc;
                end
                211: begin
                        tc = f210;
                        p32 = p32 - tc;
                        p195 = p195 + tc;
                        p213 = p213 + tc;
                end
                212: begin
                        tc = f211;
                        p213 = p213 - tc;
                        p32 = p32 + tc;
                end
                213: begin
                        tc = f212;
                        p215 = p215 - tc;
                        p214 = p214 + tc;
                end
                214: begin
                        tc = f213;
                        p216 = p216 - tc;
                        p215 = p215 + tc;
                end
                215: begin
                        tc = f214;
                        p210 = p210 - tc;
                        p214 = p214 - tc;
                        p25 = p25 + tc;
                end
                216: begin
                        tc = f215;
                        p196 = p196 - tc;
                        p212 = p212 + tc;
                        p216 = p216 + tc;
                end
                217: begin
                        tc = f216;
                        p197 = p197 - tc;
                        p33 = p33 + tc;
                end
                218: begin
                        tc = f217;
                        p33 = p33 - tc;
                end
                219: begin
                        tc = f218;
                        p217 = p217 - tc;
                        p198 = p198 + tc;
                end
                220: begin
                        tc = f219;
                        p26 = p26 - tc;
                        p217 = p217 + tc;
                end
                221: begin
                        tc = f220;
                        p219 = p219 - tc;
                        p220 = p220 + tc;
                end
                222: begin
                        tc = f221;
                        p222 = p222 - tc;
                        p221 = p221 + tc;
                end
                223: begin
                        tc = f222;
                        p30 = p30 - tc;
                        p218 = p218 + tc;
                        p223 = p223 + tc;
                end
                224: begin
                        tc = f223;
                        p223 = p223 - tc;
                        p30 = p30 + tc;
                end
                225: begin
                        tc = f224;
                        p225 = p225 - tc;
                        p224 = p224 + tc;
                end
                226: begin
                        tc = f225;
                        p226 = p226 - tc;
                        p225 = p225 + tc;
                end
                227: begin
                        tc = f226;
                        p33 = p33 - tc;
                        p219 = p219 + tc;
                        p227 = p227 + tc;
                end
                228: begin
                        tc = f227;
                        p227 = p227 - tc;
                        p33 = p33 + tc;
                end
                229: begin
                        tc = f228;
                        p229 = p229 - tc;
                        p228 = p228 + tc;
                end
                230: begin
                        tc = f229;
                        p230 = p230 - tc;
                        p229 = p229 + tc;
                end
                231: begin
                        tc = f230;
                        p224 = p224 - tc;
                        p228 = p228 - tc;
                        p26 = p26 + tc;
                end
                232: begin
                        tc = f231;
                        p221 = p221 - tc;
                        p226 = p226 + tc;
                        p230 = p230 + tc;
                end
                233: begin
                        tc = f232;
                        p220 = p220 - tc;
                        p34 = p34 + tc;
                end
                234: begin
                        tc = f233;
                        p34 = p34 - tc;
                end
                235: begin
                        tc = f234;
                        p231 = p231 - tc;
                        p222 = p222 + tc;
                end
                236: begin
                        tc = f235;
                        p27 = p27 - tc;
                        p231 = p231 + tc;
                end
                237: begin
                        tc = f236;
                        p238 = p238 - tc;
                        p234 = p234 + tc;
                end
                238: begin
                        tc = f237;
                        p232 = p232 - tc;
                end
                239: begin
                        tc = f238;
                        p236 = p236 - tc;
                        p238 = p238 + tc;
                end
                240: begin
                        tc = f239;
                        p233 = p233 - tc*2;
                        p239 = p239 + tc;
                end
                241: begin
                        tc = f240;
                        p240 = p240 - tc;
                        p237 = p237 + tc;
                end
                242: begin
                        tc = f241;
                        p233 = p233 - tc;
                        p242 = p242 - tc;
                        p241 = p241 + tc;
                end
                243: begin
                        tc = f242;
                        p243 = p243 - tc;
                        p240 = p240 + tc;
                end
                244: begin
                        tc = f243;
                        p232 = p232 - tc;
                        p235 = p235 + tc;
                        p244 = p244 + tc;
                end
                245: begin
                        tc = f244;
                        p232 = p232 - tc;
                        p244 = p244 + tc;
                end
                246: begin
                        tc = f245;
                        p245 = p245 - tc;
                        p243 = p243 + tc;
                end
                247: begin
                        tc = f246;
                        p239 = p239 - tc;
                        p233 = p233 + tc;
                end
                248: begin
                        tc = f247;
                        p246 = p246 - tc;
                        p245 = p245 + tc;
                end
                249: begin
                        tc = f248;
                        p244 = p244 - tc;
                        p232 = p232 + tc*2;
                end
                250: begin
                        tc = f249;
                        p234 = p234 - tc;
                        p241 = p241 - tc;
                        p242 = p242 + tc;
                        p246 = p246 + tc;
                end
                251: begin
                        tc = f250;
                        p234 = p234 - tc;
                        p246 = p246 + tc;
                end
                252: begin
                        tc = f251;
                        p39 = p39 - tc;
                        p232 = p232 + tc;
                        p247 = p247 + tc;
                end
                253: begin
                        tc = f252;
                        p247 = p247 - tc;
                        p39 = p39 + tc;
                end
                254: begin
                        tc = f253;
                        p249 = p249 - tc;
                        p248 = p248 + tc;
                end
                255: begin
                        tc = f254;
                        p250 = p250 - tc;
                        p249 = p249 + tc;
                end
                256: begin
                        tc = f255;
                        p40 = p40 - tc;
                        p233 = p233 + tc;
                        p251 = p251 + tc;
                end
                257: begin
                        tc = f256;
                        p251 = p251 - tc;
                        p40 = p40 + tc;
                end
                258: begin
                        tc = f257;
                        p253 = p253 - tc;
                        p252 = p252 + tc;
                end
                259: begin
                        tc = f258;
                        p254 = p254 - tc;
                        p253 = p253 + tc;
                end
                260: begin
                        tc = f259;
                        p248 = p248 - tc;
                        p252 = p252 - tc;
                        p35 = p35 + tc;
                end
                261: begin
                        tc = f260;
                        p234 = p234 - tc;
                        p250 = p250 + tc;
                        p254 = p254 + tc;
                end
                262: begin
                        tc = f261;
                        p235 = p235 - tc;
                        p41 = p41 + tc;
                end
                263: begin
                        tc = f262;
                        p41 = p41 - tc;
                end
                264: begin
                        tc = f263;
                        p255 = p255 - tc;
                        p236 = p236 + tc;
                end
                265: begin
                        tc = f264;
                        p36 = p36 - tc;
                        p255 = p255 + tc;
                end
                266: begin
                        tc = f265;
                        p262 = p262 - tc;
                        p258 = p258 + tc;
                end
                267: begin
                        tc = f266;
                        p256 = p256 - tc;
                end
                268: begin
                        tc = f267;
                        p260 = p260 - tc;
                        p262 = p262 + tc;
                end
                269: begin
                        tc = f268;
                        p257 = p257 - tc*2;
                        p263 = p263 + tc;
                end
                270: begin
                        tc = f269;
                        p264 = p264 - tc;
                        p261 = p261 + tc;
                end
                271: begin
                        tc = f270;
                        p257 = p257 - tc;
                        p266 = p266 - tc;
                        p265 = p265 + tc;
                end
                272: begin
                        tc = f271;
                        p267 = p267 - tc;
                        p264 = p264 + tc;
                end
                273: begin
                        tc = f272;
                        p256 = p256 - tc;
                        p259 = p259 + tc;
                        p268 = p268 + tc;
                end
                274: begin
                        tc = f273;
                        p256 = p256 - tc;
                        p268 = p268 + tc;
                end
                275: begin
                        tc = f274;
                        p269 = p269 - tc;
                        p267 = p267 + tc;
                end
                276: begin
                        tc = f275;
                        p263 = p263 - tc;
                        p257 = p257 + tc;
                end
                277: begin
                        tc = f276;
                        p270 = p270 - tc;
                        p269 = p269 + tc;
                end
                278: begin
                        tc = f277;
                        p268 = p268 - tc;
                        p256 = p256 + tc*2;
                end
                279: begin
                        tc = f278;
                        p258 = p258 - tc;
                        p265 = p265 - tc;
                        p266 = p266 + tc;
                        p270 = p270 + tc;
                end
                280: begin
                        tc = f279;
                        p258 = p258 - tc;
                        p270 = p270 + tc;
                end
                281: begin
                        tc = f280;
                        p42 = p42 - tc;
                        p256 = p256 + tc;
                        p271 = p271 + tc;
                end
                282: begin
                        tc = f281;
                        p271 = p271 - tc;
                        p42 = p42 + tc;
                end
                283: begin
                        tc = f282;
                        p273 = p273 - tc;
                        p272 = p272 + tc;
                end
                284: begin
                        tc = f283;
                        p274 = p274 - tc;
                        p273 = p273 + tc;
                end
                285: begin
                        tc = f284;
                        p43 = p43 - tc;
                        p257 = p257 + tc;
                        p275 = p275 + tc;
                end
                286: begin
                        tc = f285;
                        p275 = p275 - tc;
                        p43 = p43 + tc;
                end
                287: begin
                        tc = f286;
                        p277 = p277 - tc;
                        p276 = p276 + tc;
                end
                288: begin
                        tc = f287;
                        p278 = p278 - tc;
                        p277 = p277 + tc;
                end
                289: begin
                        tc = f288;
                        p272 = p272 - tc;
                        p276 = p276 - tc;
                        p36 = p36 + tc;
                end
                290: begin
                        tc = f289;
                        p258 = p258 - tc;
                        p274 = p274 + tc;
                        p278 = p278 + tc;
                end
                291: begin
                        tc = f290;
                        p259 = p259 - tc;
                        p44 = p44 + tc;
                end
                292: begin
                        tc = f291;
                        p44 = p44 - tc;
                end
                293: begin
                        tc = f292;
                        p279 = p279 - tc;
                        p260 = p260 + tc;
                end
                294: begin
                        tc = f293;
                        p37 = p37 - tc;
                        p279 = p279 + tc;
                end
                295: begin
                        tc = f294;
                        p281 = p281 - tc;
                        p282 = p282 + tc;
                end
                296: begin
                        tc = f295;
                        p284 = p284 - tc;
                        p283 = p283 + tc;
                end
                297: begin
                        tc = f296;
                        p41 = p41 - tc;
                        p280 = p280 + tc;
                        p285 = p285 + tc;
                end
                298: begin
                        tc = f297;
                        p285 = p285 - tc;
                        p41 = p41 + tc;
                end
                299: begin
                        tc = f298;
                        p287 = p287 - tc;
                        p286 = p286 + tc;
                end
                300: begin
                        tc = f299;
                        p288 = p288 - tc;
                        p287 = p287 + tc;
                end
                301: begin
                        tc = f300;
                        p44 = p44 - tc;
                        p281 = p281 + tc;
                        p289 = p289 + tc;
                end
                302: begin
                        tc = f301;
                        p289 = p289 - tc;
                        p44 = p44 + tc;
                end
                303: begin
                        tc = f302;
                        p291 = p291 - tc;
                        p290 = p290 + tc;
                end
                304: begin
                        tc = f303;
                        p292 = p292 - tc;
                        p291 = p291 + tc;
                end
                305: begin
                        tc = f304;
                        p286 = p286 - tc;
                        p290 = p290 - tc;
                        p37 = p37 + tc;
                end
                306: begin
                        tc = f305;
                        p283 = p283 - tc;
                        p288 = p288 + tc;
                        p292 = p292 + tc;
                end
                307: begin
                        tc = f306;
                        p282 = p282 - tc;
                        p45 = p45 + tc;
                end
                308: begin
                        tc = f307;
                        p45 = p45 - tc;
                end
                309: begin
                        tc = f308;
                        p293 = p293 - tc;
                        p284 = p284 + tc;
                end
                310: begin
                        tc = f309;
                        p38 = p38 - tc;
                        p293 = p293 + tc;
                end
                default:;
        endcase
//        led = ~p12[5:0];
        if(tf>0) counter1=counter1+1;
end
end
reg [32:0] counter;

always @(posedge clk) begin
    if (counter < 32'd2_7500_0000)       //delay
        counter <= counter + 1'b1;
    else
        counter <= 32'd0;
end

always @(posedge clk) begin
    if (counter == 32'd0)       
        led <= ~counter1[47:42];
    else if (counter == 32'd2500_0000)       
        led <= ~counter1[41:36];
    else if (counter == 32'd5000_0000)       
        led <= ~counter1[35:30];
    else if (counter == 32'd7500_0000)       
        led <= ~counter1[29:24];
    else if (counter == 32'd1_0000_0000)       
        led <= ~counter1[23:18];
    else if (counter == 32'd1_2500_0000)       
        led <= ~counter1[17:12];
    else if (counter == 32'd1_5000_0000)       
        led <= ~counter1[11:6];
    else if (counter == 32'd1_7500_0000)       
        led <= ~counter1[5:0];
    else if (counter == 32'd2_0000_0000)       
        led <= 6'b000000;
    else if (counter == 32'd2_2500_0000)       
        led <= 6'b111111;
    else if (counter == 32'd2_5000_0000)       
        led <= 6'b000000;
    else
        led <= led;
end
endmodule