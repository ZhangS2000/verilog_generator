module sn(
        input clk,
        output reg [5:0] led
);
`define INH(place) ((place) == 0 ? 131071 : 0)
reg [16:0] p0=0,p1=1,p2=1,p3=1,p4=1,p5=1,p6=1,p7=1,p8=1,p9=1,p10=8,p11=20,p12=0,p13=20,p14=0,p15=20,p16=0,p17=5,p18=20,p19=0,p20=20,p21=0,p22=0,p23=1,p24=20,p25=0,p26=0,p27=10,p28=0,p29=0,p30=0,p31=1,p32=0,p33=1,p34=1,p35=1,p36=0,p37=1,p38=0,p39=1,p40=1,p41=0,p42=1,p43=1,p44=0,p45=1,p46=1,p47=1,p48=0,p49=1,p50=1,p51=1,p52=1,p53=0,p54=0,p55=1,p56=0,p57=1,p58=1,p59=1,p60=0,p61=1,p62=0,p63=1,p64=1,p65=0,p66=1,p67=1,p68=0,p69=1,p70=1,p71=1,p72=0,p73=1,p74=1,p75=1,p76=1,p77=0,p78=0,p79=1,p80=0,p81=1,p82=1,p83=1,p84=0,p85=1,p86=0,p87=1,p88=1,p89=0,p90=1,p91=1,p92=0,p93=1,p94=1,p95=1,p96=0,p97=1,p98=1,p99=1,p100=1,p101=0,p102=0,p103=1,p104=0,p105=1,p106=1,p107=1,p108=0,p109=1,p110=0,p111=1,p112=1,p113=0,p114=1,p115=1,p116=0,p117=1,p118=1,p119=1,p120=0,p121=1,p122=1,p123=1,p124=1,p125=0,p126=0,p127=1,p128=0,p129=1,p130=1,p131=1,p132=0,p133=1,p134=0,p135=1,p136=1,p137=0,p138=1,p139=1,p140=0,p141=1,p142=1,p143=1,p144=0,p145=1,p146=1,p147=1,p148=1,p149=0,p150=0,p151=0,p152=1,p153=1,p154=0,p155=1,p156=1,p157=1,p158=0,p159=1,p160=1,p161=1,p162=1,p163=0,p164=0,p165=1,p166=0,p167=1,p168=1,p169=1,p170=0,p171=1,p172=0,p173=1,p174=1,p175=0,p176=1,p177=1,p178=0,p179=1,p180=1,p181=1,p182=0,p183=1,p184=1,p185=1,p186=1,p187=0,p188=0,p189=0,p190=1,p191=1,p192=0,p193=1,p194=1,p195=1,p196=0,p197=1,p198=1,p199=1,p200=1,p201=0,p202=0,p203=0,p204=1,p205=1,p206=0,p207=1,p208=1,p209=1,p210=0,p211=1,p212=1,p213=1,p214=1;
reg [16:0] f0,f1,f2,f3,f4,f5,f6,f7,f8,f9,f10,f11,f12,f13,f14,f15,f16,f17,f18,f19,f20,f21,f22,f23,f24,f25,f26,f27,f28,f29,f30,f31,f32,f33,f34,f35,f36,f37,f38,f39,f40,f41,f42,f43,f44,f45,f46,f47,f48,f49,f50,f51,f52,f53,f54,f55,f56,f57,f58,f59,f60,f61,f62,f63,f64,f65,f66,f67,f68,f69,f70,f71,f72,f73,f74,f75,f76,f77,f78,f79,f80,f81,f82,f83,f84,f85,f86,f87,f88,f89,f90,f91,f92,f93,f94,f95,f96,f97,f98,f99,f100,f101,f102,f103,f104,f105,f106,f107,f108,f109,f110,f111,f112,f113,f114,f115,f116,f117,f118,f119,f120,f121,f122,f123,f124,f125,f126,f127,f128,f129,f130,f131,f132,f133,f134,f135,f136,f137,f138,f139,f140,f141,f142,f143,f144,f145,f146,f147,f148,f149,f150,f151,f152,f153,f154,f155,f156,f157,f158,f159,f160,f161,f162,f163,f164,f165,f166,f167,f168,f169,f170,f171,f172,f173,f174,f175,f176,f177,f178,f179,f180,f181,f182,f183,f184,f185,f186,f187,f188,f189,f190,f191,f192,f193,f194,f195,f196,f197,f198,f199,f200,f201,f202,f203,f204,f205,f206,f207,f208,f209,f210,f211,f212,f213,f214,f215,f216,f217,f218,f219,f220,f221,f222,f223,f224,f225,f226,f227,f228,f229,f230;
reg [16:0] tf;
reg [16:0] tc;
reg [47:0] counter1=1;
reg [1:0] clk_div; // 2位寄存器用于实现时钟分频

always @(posedge clk) begin
    if(clk_div < 2'b01)
        clk_div <= clk_div + 1; // 计数器自增
    else
        clk_div <= 2'b00; // 重置计数器
end

// 使用clk_div来控制某些逻辑的触发条件
always @(posedge clk) begin
    if (clk_div == 2'b01) begin
        f0 = 131071;
        f0 = (f0 >= `INH(p31)) ? `INH(p31) : f0;
        f0 = (f0 > p34) ? p34 : f0;
        f1 = 131071;
        f1 = (f1 >= `INH(p55)) ? `INH(p55) : f1;
        f1 = (f1 > p58) ? p58 : f1;
        f2 = 131071;
        f2 = (f2 >= `INH(p79)) ? `INH(p79) : f2;
        f2 = (f2 > p82) ? p82 : f2;
        f3 = 131071;
        f3 = (f3 >= `INH(p103)) ? `INH(p103) : f3;
        f3 = (f3 > p106) ? p106 : f3;
        f4 = 131071;
        f4 = (f4 >= `INH(p127)) ? `INH(p127) : f4;
        f4 = (f4 > p130) ? p130 : f4;
        f5 = 131071;
        f5 = (f5 > p149) ? p149 : f5;
        f5 = (f5 >= `INH(p152)) ? `INH(p152) : f5;
        f6 = 131071;
        f6 = (f6 >= `INH(p165)) ? `INH(p165) : f6;
        f6 = (f6 > p168) ? p168 : f6;
        f7 = 131071;
        f7 = (f7 > p187) ? p187 : f7;
        f7 = (f7 >= `INH(p190)) ? `INH(p190) : f7;
        f8 = 131071;
        f8 = (f8 > p201) ? p201 : f8;
        f8 = (f8 >= `INH(p204)) ? `INH(p204) : f8;
        f9 = 131071;
        f9 = (f9 >= `INH(p30)) ? `INH(p30) : f9;
        f9 = (f9 >= `INH(p31)) ? `INH(p31) : f9;
        f9 = (f9 > p35) ? p35 : f9;
        f10 = 131071;
        f10 = (f10 > p29) ? p29 : f10;
        f10 = (f10 >= `INH(p35)) ? `INH(p35) : f10;
        f11 = 131071;
        f11 = (f11 > p33) ? p33 : f11;
        f11 = (f11 >= `INH(p35)) ? `INH(p35) : f11;
        f12 = 131071;
        f12 = (f12 >= p30/2) ? p30/2 : f12;
        f12 = (f12 >= `INH(p34)) ? `INH(p34) : f12;
        f13 = 131071;
        f13 = (f13 >= `INH(p34)) ? `INH(p34) : f13;
        f13 = (f13 > p37) ? p37 : f13;
        f14 = 131071;
        f14 = (f14 > p30) ? p30 : f14;
        f14 = (f14 >= `INH(p37)) ? `INH(p37) : f14;
        f14 = (f14 > p39) ? p39 : f14;
        f15 = 131071;
        f15 = (f15 >= `INH(p37)) ? `INH(p37) : f15;
        f15 = (f15 > p40) ? p40 : f15;
        f16 = 131071;
        f16 = (f16 > p29) ? p29 : f16;
        f16 = (f16 >= `INH(p39)) ? `INH(p39) : f16;
        f16 = (f16 >= `INH(p40)) ? `INH(p40) : f16;
        f17 = 131071;
        f17 = (f17 > p29) ? p29 : f17;
        f17 = (f17 >= `INH(p38)) ? `INH(p38) : f17;
        f17 = (f17 >= `INH(p40)) ? `INH(p40) : f17;
        f18 = 131071;
        f18 = (f18 >= `INH(p40)) ? `INH(p40) : f18;
        f18 = (f18 > p42) ? p42 : f18;
        f19 = 131071;
        f19 = (f19 > p36) ? p36 : f19;
        f19 = (f19 >= `INH(p42)) ? `INH(p42) : f19;
        f20 = 131071;
        f20 = (f20 >= `INH(p42)) ? `INH(p42) : f20;
        f20 = (f20 > p43) ? p43 : f20;
        f21 = 131071;
        f21 = (f21 > p41) ? p41 : f21;
        f21 = (f21 >= `INH(p43)) ? `INH(p43) : f21;
        f22 = 131071;
        f22 = (f22 > p31) ? p31 : f22;
        f22 = (f22 > p38) ? p38 : f22;
        f22 = (f22 >= `INH(p39)) ? `INH(p39) : f22;
        f22 = (f22 >= `INH(p43)) ? `INH(p43) : f22;
        f23 = 131071;
        f23 = (f23 > p31) ? p31 : f23;
        f23 = (f23 >= `INH(p38)) ? `INH(p38) : f23;
        f23 = (f23 >= `INH(p43)) ? `INH(p43) : f23;
        f24 = 131071;
        f24 = (f24 > p10) ? p10 : f24;
        f24 = (f24 >= `INH(p45)) ? `INH(p45) : f24;
        f25 = 131071;
        f25 = (f25 > p44) ? p44 : f25;
        f25 = (f25 >= `INH(p46)) ? `INH(p46) : f25;
        f26 = 131071;
        f26 = (f26 >= `INH(p10)) ? `INH(p10) : f26;
        f26 = (f26 >= `INH(p45)) ? `INH(p45) : f26;
        f26 = (f26 > p46) ? p46 : f26;
        f27 = 131071;
        f27 = (f27 >= `INH(p44)) ? `INH(p44) : f27;
        f27 = (f27 >= `INH(p46)) ? `INH(p46) : f27;
        f27 = (f27 > p47) ? p47 : f27;
        f28 = 131071;
        f28 = (f28 > p11) ? p11 : f28;
        f28 = (f28 >= `INH(p49)) ? `INH(p49) : f28;
        f29 = 131071;
        f29 = (f29 > p48) ? p48 : f29;
        f29 = (f29 >= `INH(p50)) ? `INH(p50) : f29;
        f30 = 131071;
        f30 = (f30 >= `INH(p11)) ? `INH(p11) : f30;
        f30 = (f30 >= `INH(p49)) ? `INH(p49) : f30;
        f30 = (f30 > p50) ? p50 : f30;
        f31 = 131071;
        f31 = (f31 >= `INH(p48)) ? `INH(p48) : f31;
        f31 = (f31 >= `INH(p50)) ? `INH(p50) : f31;
        f31 = (f31 > p51) ? p51 : f31;
        f32 = 131071;
        f32 = (f32 >= `INH(p0)) ? `INH(p0) : f32;
        f32 = (f32 > p45) ? p45 : f32;
        f32 = (f32 > p49) ? p49 : f32;
        f33 = 131071;
        f33 = (f33 > p31) ? p31 : f33;
        f33 = (f33 >= `INH(p47)) ? `INH(p47) : f33;
        f33 = (f33 >= `INH(p51)) ? `INH(p51) : f33;
        f34 = 131071;
        f34 = (f34 > p32) ? p32 : f34;
        f34 = (f34 >= `INH(p52)) ? `INH(p52) : f34;
        f35 = 131071;
        f35 = (f35 > p12) ? p12 : f35;
        f35 = (f35 >= `INH(p33)) ? `INH(p33) : f35;
        f36 = 131071;
        f36 = (f36 >= `INH(p12)) ? `INH(p12) : f36;
        f36 = (f36 >= `INH(p33)) ? `INH(p33) : f36;
        f36 = (f36 > p52) ? p52 : f36;
        f37 = 131071;
        f37 = (f37 > p1) ? p1 : f37;
        f37 = (f37 >= `INH(p32)) ? `INH(p32) : f37;
        f37 = (f37 >= `INH(p52)) ? `INH(p52) : f37;
        f38 = 131071;
        f38 = (f38 >= `INH(p54)) ? `INH(p54) : f38;
        f38 = (f38 >= `INH(p55)) ? `INH(p55) : f38;
        f38 = (f38 > p59) ? p59 : f38;
        f39 = 131071;
        f39 = (f39 > p53) ? p53 : f39;
        f39 = (f39 >= `INH(p59)) ? `INH(p59) : f39;
        f40 = 131071;
        f40 = (f40 > p57) ? p57 : f40;
        f40 = (f40 >= `INH(p59)) ? `INH(p59) : f40;
        f41 = 131071;
        f41 = (f41 >= p54/2) ? p54/2 : f41;
        f41 = (f41 >= `INH(p58)) ? `INH(p58) : f41;
        f42 = 131071;
        f42 = (f42 >= `INH(p58)) ? `INH(p58) : f42;
        f42 = (f42 > p61) ? p61 : f42;
        f43 = 131071;
        f43 = (f43 > p54) ? p54 : f43;
        f43 = (f43 >= `INH(p61)) ? `INH(p61) : f43;
        f43 = (f43 > p63) ? p63 : f43;
        f44 = 131071;
        f44 = (f44 >= `INH(p61)) ? `INH(p61) : f44;
        f44 = (f44 > p64) ? p64 : f44;
        f45 = 131071;
        f45 = (f45 > p53) ? p53 : f45;
        f45 = (f45 >= `INH(p63)) ? `INH(p63) : f45;
        f45 = (f45 >= `INH(p64)) ? `INH(p64) : f45;
        f46 = 131071;
        f46 = (f46 > p53) ? p53 : f46;
        f46 = (f46 >= `INH(p62)) ? `INH(p62) : f46;
        f46 = (f46 >= `INH(p64)) ? `INH(p64) : f46;
        f47 = 131071;
        f47 = (f47 >= `INH(p64)) ? `INH(p64) : f47;
        f47 = (f47 > p66) ? p66 : f47;
        f48 = 131071;
        f48 = (f48 > p60) ? p60 : f48;
        f48 = (f48 >= `INH(p66)) ? `INH(p66) : f48;
        f49 = 131071;
        f49 = (f49 >= `INH(p66)) ? `INH(p66) : f49;
        f49 = (f49 > p67) ? p67 : f49;
        f50 = 131071;
        f50 = (f50 > p65) ? p65 : f50;
        f50 = (f50 >= `INH(p67)) ? `INH(p67) : f50;
        f51 = 131071;
        f51 = (f51 > p55) ? p55 : f51;
        f51 = (f51 > p62) ? p62 : f51;
        f51 = (f51 >= `INH(p63)) ? `INH(p63) : f51;
        f51 = (f51 >= `INH(p67)) ? `INH(p67) : f51;
        f52 = 131071;
        f52 = (f52 > p55) ? p55 : f52;
        f52 = (f52 >= `INH(p62)) ? `INH(p62) : f52;
        f52 = (f52 >= `INH(p67)) ? `INH(p67) : f52;
        f53 = 131071;
        f53 = (f53 > p12) ? p12 : f53;
        f53 = (f53 >= `INH(p69)) ? `INH(p69) : f53;
        f54 = 131071;
        f54 = (f54 > p68) ? p68 : f54;
        f54 = (f54 >= `INH(p70)) ? `INH(p70) : f54;
        f55 = 131071;
        f55 = (f55 >= `INH(p12)) ? `INH(p12) : f55;
        f55 = (f55 >= `INH(p69)) ? `INH(p69) : f55;
        f55 = (f55 > p70) ? p70 : f55;
        f56 = 131071;
        f56 = (f56 >= `INH(p68)) ? `INH(p68) : f56;
        f56 = (f56 >= `INH(p70)) ? `INH(p70) : f56;
        f56 = (f56 > p71) ? p71 : f56;
        f57 = 131071;
        f57 = (f57 > p13) ? p13 : f57;
        f57 = (f57 >= `INH(p73)) ? `INH(p73) : f57;
        f58 = 131071;
        f58 = (f58 > p72) ? p72 : f58;
        f58 = (f58 >= `INH(p74)) ? `INH(p74) : f58;
        f59 = 131071;
        f59 = (f59 >= `INH(p13)) ? `INH(p13) : f59;
        f59 = (f59 >= `INH(p73)) ? `INH(p73) : f59;
        f59 = (f59 > p74) ? p74 : f59;
        f60 = 131071;
        f60 = (f60 >= `INH(p72)) ? `INH(p72) : f60;
        f60 = (f60 >= `INH(p74)) ? `INH(p74) : f60;
        f60 = (f60 > p75) ? p75 : f60;
        f61 = 131071;
        f61 = (f61 >= `INH(p1)) ? `INH(p1) : f61;
        f61 = (f61 > p69) ? p69 : f61;
        f61 = (f61 > p73) ? p73 : f61;
        f62 = 131071;
        f62 = (f62 > p55) ? p55 : f62;
        f62 = (f62 >= `INH(p71)) ? `INH(p71) : f62;
        f62 = (f62 >= `INH(p75)) ? `INH(p75) : f62;
        f63 = 131071;
        f63 = (f63 > p56) ? p56 : f63;
        f63 = (f63 >= `INH(p76)) ? `INH(p76) : f63;
        f64 = 131071;
        f64 = (f64 > p14) ? p14 : f64;
        f64 = (f64 >= `INH(p57)) ? `INH(p57) : f64;
        f65 = 131071;
        f65 = (f65 >= `INH(p14)) ? `INH(p14) : f65;
        f65 = (f65 >= `INH(p57)) ? `INH(p57) : f65;
        f65 = (f65 > p76) ? p76 : f65;
        f66 = 131071;
        f66 = (f66 > p2) ? p2 : f66;
        f66 = (f66 >= `INH(p56)) ? `INH(p56) : f66;
        f66 = (f66 >= `INH(p76)) ? `INH(p76) : f66;
        f67 = 131071;
        f67 = (f67 >= `INH(p78)) ? `INH(p78) : f67;
        f67 = (f67 >= `INH(p79)) ? `INH(p79) : f67;
        f67 = (f67 > p83) ? p83 : f67;
        f68 = 131071;
        f68 = (f68 > p77) ? p77 : f68;
        f68 = (f68 >= `INH(p83)) ? `INH(p83) : f68;
        f69 = 131071;
        f69 = (f69 > p81) ? p81 : f69;
        f69 = (f69 >= `INH(p83)) ? `INH(p83) : f69;
        f70 = 131071;
        f70 = (f70 >= p78/2) ? p78/2 : f70;
        f70 = (f70 >= `INH(p82)) ? `INH(p82) : f70;
        f71 = 131071;
        f71 = (f71 >= `INH(p82)) ? `INH(p82) : f71;
        f71 = (f71 > p85) ? p85 : f71;
        f72 = 131071;
        f72 = (f72 > p78) ? p78 : f72;
        f72 = (f72 >= `INH(p85)) ? `INH(p85) : f72;
        f72 = (f72 > p87) ? p87 : f72;
        f73 = 131071;
        f73 = (f73 >= `INH(p85)) ? `INH(p85) : f73;
        f73 = (f73 > p88) ? p88 : f73;
        f74 = 131071;
        f74 = (f74 > p77) ? p77 : f74;
        f74 = (f74 >= `INH(p87)) ? `INH(p87) : f74;
        f74 = (f74 >= `INH(p88)) ? `INH(p88) : f74;
        f75 = 131071;
        f75 = (f75 > p77) ? p77 : f75;
        f75 = (f75 >= `INH(p86)) ? `INH(p86) : f75;
        f75 = (f75 >= `INH(p88)) ? `INH(p88) : f75;
        f76 = 131071;
        f76 = (f76 >= `INH(p88)) ? `INH(p88) : f76;
        f76 = (f76 > p90) ? p90 : f76;
        f77 = 131071;
        f77 = (f77 > p84) ? p84 : f77;
        f77 = (f77 >= `INH(p90)) ? `INH(p90) : f77;
        f78 = 131071;
        f78 = (f78 >= `INH(p90)) ? `INH(p90) : f78;
        f78 = (f78 > p91) ? p91 : f78;
        f79 = 131071;
        f79 = (f79 > p89) ? p89 : f79;
        f79 = (f79 >= `INH(p91)) ? `INH(p91) : f79;
        f80 = 131071;
        f80 = (f80 > p79) ? p79 : f80;
        f80 = (f80 > p86) ? p86 : f80;
        f80 = (f80 >= `INH(p87)) ? `INH(p87) : f80;
        f80 = (f80 >= `INH(p91)) ? `INH(p91) : f80;
        f81 = 131071;
        f81 = (f81 > p79) ? p79 : f81;
        f81 = (f81 >= `INH(p86)) ? `INH(p86) : f81;
        f81 = (f81 >= `INH(p91)) ? `INH(p91) : f81;
        f82 = 131071;
        f82 = (f82 > p14) ? p14 : f82;
        f82 = (f82 >= `INH(p93)) ? `INH(p93) : f82;
        f83 = 131071;
        f83 = (f83 > p92) ? p92 : f83;
        f83 = (f83 >= `INH(p94)) ? `INH(p94) : f83;
        f84 = 131071;
        f84 = (f84 >= `INH(p14)) ? `INH(p14) : f84;
        f84 = (f84 >= `INH(p93)) ? `INH(p93) : f84;
        f84 = (f84 > p94) ? p94 : f84;
        f85 = 131071;
        f85 = (f85 >= `INH(p92)) ? `INH(p92) : f85;
        f85 = (f85 >= `INH(p94)) ? `INH(p94) : f85;
        f85 = (f85 > p95) ? p95 : f85;
        f86 = 131071;
        f86 = (f86 > p15) ? p15 : f86;
        f86 = (f86 >= `INH(p97)) ? `INH(p97) : f86;
        f87 = 131071;
        f87 = (f87 > p96) ? p96 : f87;
        f87 = (f87 >= `INH(p98)) ? `INH(p98) : f87;
        f88 = 131071;
        f88 = (f88 >= `INH(p15)) ? `INH(p15) : f88;
        f88 = (f88 >= `INH(p97)) ? `INH(p97) : f88;
        f88 = (f88 > p98) ? p98 : f88;
        f89 = 131071;
        f89 = (f89 >= `INH(p96)) ? `INH(p96) : f89;
        f89 = (f89 >= `INH(p98)) ? `INH(p98) : f89;
        f89 = (f89 > p99) ? p99 : f89;
        f90 = 131071;
        f90 = (f90 >= `INH(p2)) ? `INH(p2) : f90;
        f90 = (f90 > p93) ? p93 : f90;
        f90 = (f90 > p97) ? p97 : f90;
        f91 = 131071;
        f91 = (f91 > p79) ? p79 : f91;
        f91 = (f91 >= `INH(p95)) ? `INH(p95) : f91;
        f91 = (f91 >= `INH(p99)) ? `INH(p99) : f91;
        f92 = 131071;
        f92 = (f92 > p80) ? p80 : f92;
        f92 = (f92 >= `INH(p100)) ? `INH(p100) : f92;
        f93 = 131071;
        f93 = (f93 > p16) ? p16 : f93;
        f93 = (f93 >= `INH(p81)) ? `INH(p81) : f93;
        f94 = 131071;
        f94 = (f94 >= `INH(p16)) ? `INH(p16) : f94;
        f94 = (f94 >= `INH(p81)) ? `INH(p81) : f94;
        f94 = (f94 > p100) ? p100 : f94;
        f95 = 131071;
        f95 = (f95 > p3) ? p3 : f95;
        f95 = (f95 >= `INH(p80)) ? `INH(p80) : f95;
        f95 = (f95 >= `INH(p100)) ? `INH(p100) : f95;
        f96 = 131071;
        f96 = (f96 >= `INH(p102)) ? `INH(p102) : f96;
        f96 = (f96 >= `INH(p103)) ? `INH(p103) : f96;
        f96 = (f96 > p107) ? p107 : f96;
        f97 = 131071;
        f97 = (f97 > p101) ? p101 : f97;
        f97 = (f97 >= `INH(p107)) ? `INH(p107) : f97;
        f98 = 131071;
        f98 = (f98 > p105) ? p105 : f98;
        f98 = (f98 >= `INH(p107)) ? `INH(p107) : f98;
        f99 = 131071;
        f99 = (f99 >= p102/2) ? p102/2 : f99;
        f99 = (f99 >= `INH(p106)) ? `INH(p106) : f99;
        f100 = 131071;
        f100 = (f100 >= `INH(p106)) ? `INH(p106) : f100;
        f100 = (f100 > p109) ? p109 : f100;
        f101 = 131071;
        f101 = (f101 > p102) ? p102 : f101;
        f101 = (f101 >= `INH(p109)) ? `INH(p109) : f101;
        f101 = (f101 > p111) ? p111 : f101;
        f102 = 131071;
        f102 = (f102 >= `INH(p109)) ? `INH(p109) : f102;
        f102 = (f102 > p112) ? p112 : f102;
        f103 = 131071;
        f103 = (f103 > p101) ? p101 : f103;
        f103 = (f103 >= `INH(p111)) ? `INH(p111) : f103;
        f103 = (f103 >= `INH(p112)) ? `INH(p112) : f103;
        f104 = 131071;
        f104 = (f104 > p101) ? p101 : f104;
        f104 = (f104 >= `INH(p110)) ? `INH(p110) : f104;
        f104 = (f104 >= `INH(p112)) ? `INH(p112) : f104;
        f105 = 131071;
        f105 = (f105 >= `INH(p112)) ? `INH(p112) : f105;
        f105 = (f105 > p114) ? p114 : f105;
        f106 = 131071;
        f106 = (f106 > p108) ? p108 : f106;
        f106 = (f106 >= `INH(p114)) ? `INH(p114) : f106;
        f107 = 131071;
        f107 = (f107 >= `INH(p114)) ? `INH(p114) : f107;
        f107 = (f107 > p115) ? p115 : f107;
        f108 = 131071;
        f108 = (f108 > p113) ? p113 : f108;
        f108 = (f108 >= `INH(p115)) ? `INH(p115) : f108;
        f109 = 131071;
        f109 = (f109 > p103) ? p103 : f109;
        f109 = (f109 > p110) ? p110 : f109;
        f109 = (f109 >= `INH(p111)) ? `INH(p111) : f109;
        f109 = (f109 >= `INH(p115)) ? `INH(p115) : f109;
        f110 = 131071;
        f110 = (f110 > p103) ? p103 : f110;
        f110 = (f110 >= `INH(p110)) ? `INH(p110) : f110;
        f110 = (f110 >= `INH(p115)) ? `INH(p115) : f110;
        f111 = 131071;
        f111 = (f111 > p17) ? p17 : f111;
        f111 = (f111 >= `INH(p117)) ? `INH(p117) : f111;
        f112 = 131071;
        f112 = (f112 > p116) ? p116 : f112;
        f112 = (f112 >= `INH(p118)) ? `INH(p118) : f112;
        f113 = 131071;
        f113 = (f113 >= `INH(p17)) ? `INH(p17) : f113;
        f113 = (f113 >= `INH(p117)) ? `INH(p117) : f113;
        f113 = (f113 > p118) ? p118 : f113;
        f114 = 131071;
        f114 = (f114 >= `INH(p116)) ? `INH(p116) : f114;
        f114 = (f114 >= `INH(p118)) ? `INH(p118) : f114;
        f114 = (f114 > p119) ? p119 : f114;
        f115 = 131071;
        f115 = (f115 > p18) ? p18 : f115;
        f115 = (f115 >= `INH(p121)) ? `INH(p121) : f115;
        f116 = 131071;
        f116 = (f116 > p120) ? p120 : f116;
        f116 = (f116 >= `INH(p122)) ? `INH(p122) : f116;
        f117 = 131071;
        f117 = (f117 >= `INH(p18)) ? `INH(p18) : f117;
        f117 = (f117 >= `INH(p121)) ? `INH(p121) : f117;
        f117 = (f117 > p122) ? p122 : f117;
        f118 = 131071;
        f118 = (f118 >= `INH(p120)) ? `INH(p120) : f118;
        f118 = (f118 >= `INH(p122)) ? `INH(p122) : f118;
        f118 = (f118 > p123) ? p123 : f118;
        f119 = 131071;
        f119 = (f119 >= `INH(p3)) ? `INH(p3) : f119;
        f119 = (f119 > p117) ? p117 : f119;
        f119 = (f119 > p121) ? p121 : f119;
        f120 = 131071;
        f120 = (f120 > p103) ? p103 : f120;
        f120 = (f120 >= `INH(p119)) ? `INH(p119) : f120;
        f120 = (f120 >= `INH(p123)) ? `INH(p123) : f120;
        f121 = 131071;
        f121 = (f121 > p104) ? p104 : f121;
        f121 = (f121 >= `INH(p124)) ? `INH(p124) : f121;
        f122 = 131071;
        f122 = (f122 > p19) ? p19 : f122;
        f122 = (f122 >= `INH(p105)) ? `INH(p105) : f122;
        f123 = 131071;
        f123 = (f123 >= `INH(p19)) ? `INH(p19) : f123;
        f123 = (f123 >= `INH(p105)) ? `INH(p105) : f123;
        f123 = (f123 > p124) ? p124 : f123;
        f124 = 131071;
        f124 = (f124 > p4) ? p4 : f124;
        f124 = (f124 >= `INH(p104)) ? `INH(p104) : f124;
        f124 = (f124 >= `INH(p124)) ? `INH(p124) : f124;
        f125 = 131071;
        f125 = (f125 >= `INH(p126)) ? `INH(p126) : f125;
        f125 = (f125 >= `INH(p127)) ? `INH(p127) : f125;
        f125 = (f125 > p131) ? p131 : f125;
        f126 = 131071;
        f126 = (f126 > p125) ? p125 : f126;
        f126 = (f126 >= `INH(p131)) ? `INH(p131) : f126;
        f127 = 131071;
        f127 = (f127 > p129) ? p129 : f127;
        f127 = (f127 >= `INH(p131)) ? `INH(p131) : f127;
        f128 = 131071;
        f128 = (f128 >= p126/2) ? p126/2 : f128;
        f128 = (f128 >= `INH(p130)) ? `INH(p130) : f128;
        f129 = 131071;
        f129 = (f129 >= `INH(p130)) ? `INH(p130) : f129;
        f129 = (f129 > p133) ? p133 : f129;
        f130 = 131071;
        f130 = (f130 > p126) ? p126 : f130;
        f130 = (f130 >= `INH(p133)) ? `INH(p133) : f130;
        f130 = (f130 > p135) ? p135 : f130;
        f131 = 131071;
        f131 = (f131 >= `INH(p133)) ? `INH(p133) : f131;
        f131 = (f131 > p136) ? p136 : f131;
        f132 = 131071;
        f132 = (f132 > p125) ? p125 : f132;
        f132 = (f132 >= `INH(p135)) ? `INH(p135) : f132;
        f132 = (f132 >= `INH(p136)) ? `INH(p136) : f132;
        f133 = 131071;
        f133 = (f133 > p125) ? p125 : f133;
        f133 = (f133 >= `INH(p134)) ? `INH(p134) : f133;
        f133 = (f133 >= `INH(p136)) ? `INH(p136) : f133;
        f134 = 131071;
        f134 = (f134 >= `INH(p136)) ? `INH(p136) : f134;
        f134 = (f134 > p138) ? p138 : f134;
        f135 = 131071;
        f135 = (f135 > p132) ? p132 : f135;
        f135 = (f135 >= `INH(p138)) ? `INH(p138) : f135;
        f136 = 131071;
        f136 = (f136 >= `INH(p138)) ? `INH(p138) : f136;
        f136 = (f136 > p139) ? p139 : f136;
        f137 = 131071;
        f137 = (f137 > p137) ? p137 : f137;
        f137 = (f137 >= `INH(p139)) ? `INH(p139) : f137;
        f138 = 131071;
        f138 = (f138 > p127) ? p127 : f138;
        f138 = (f138 > p134) ? p134 : f138;
        f138 = (f138 >= `INH(p135)) ? `INH(p135) : f138;
        f138 = (f138 >= `INH(p139)) ? `INH(p139) : f138;
        f139 = 131071;
        f139 = (f139 > p127) ? p127 : f139;
        f139 = (f139 >= `INH(p134)) ? `INH(p134) : f139;
        f139 = (f139 >= `INH(p139)) ? `INH(p139) : f139;
        f140 = 131071;
        f140 = (f140 > p19) ? p19 : f140;
        f140 = (f140 >= `INH(p141)) ? `INH(p141) : f140;
        f141 = 131071;
        f141 = (f141 > p140) ? p140 : f141;
        f141 = (f141 >= `INH(p142)) ? `INH(p142) : f141;
        f142 = 131071;
        f142 = (f142 >= `INH(p19)) ? `INH(p19) : f142;
        f142 = (f142 >= `INH(p141)) ? `INH(p141) : f142;
        f142 = (f142 > p142) ? p142 : f142;
        f143 = 131071;
        f143 = (f143 >= `INH(p140)) ? `INH(p140) : f143;
        f143 = (f143 >= `INH(p142)) ? `INH(p142) : f143;
        f143 = (f143 > p143) ? p143 : f143;
        f144 = 131071;
        f144 = (f144 > p20) ? p20 : f144;
        f144 = (f144 >= `INH(p145)) ? `INH(p145) : f144;
        f145 = 131071;
        f145 = (f145 > p144) ? p144 : f145;
        f145 = (f145 >= `INH(p146)) ? `INH(p146) : f145;
        f146 = 131071;
        f146 = (f146 >= `INH(p20)) ? `INH(p20) : f146;
        f146 = (f146 >= `INH(p145)) ? `INH(p145) : f146;
        f146 = (f146 > p146) ? p146 : f146;
        f147 = 131071;
        f147 = (f147 >= `INH(p144)) ? `INH(p144) : f147;
        f147 = (f147 >= `INH(p146)) ? `INH(p146) : f147;
        f147 = (f147 > p147) ? p147 : f147;
        f148 = 131071;
        f148 = (f148 >= `INH(p4)) ? `INH(p4) : f148;
        f148 = (f148 > p141) ? p141 : f148;
        f148 = (f148 > p145) ? p145 : f148;
        f149 = 131071;
        f149 = (f149 > p127) ? p127 : f149;
        f149 = (f149 >= `INH(p143)) ? `INH(p143) : f149;
        f149 = (f149 >= `INH(p147)) ? `INH(p147) : f149;
        f150 = 131071;
        f150 = (f150 > p128) ? p128 : f150;
        f150 = (f150 >= `INH(p148)) ? `INH(p148) : f150;
        f151 = 131071;
        f151 = (f151 > p21) ? p21 : f151;
        f151 = (f151 >= `INH(p129)) ? `INH(p129) : f151;
        f152 = 131071;
        f152 = (f152 >= `INH(p21)) ? `INH(p21) : f152;
        f152 = (f152 >= `INH(p129)) ? `INH(p129) : f152;
        f152 = (f152 > p148) ? p148 : f152;
        f153 = 131071;
        f153 = (f153 > p5) ? p5 : f153;
        f153 = (f153 >= `INH(p128)) ? `INH(p128) : f153;
        f153 = (f153 >= `INH(p148)) ? `INH(p148) : f153;
        f154 = 131071;
        f154 = (f154 > p150) ? p150 : f154;
        f154 = (f154 >= `INH(p152)) ? `INH(p152) : f154;
        f155 = 131071;
        f155 = (f155 >= `INH(p149)) ? `INH(p149) : f155;
        f155 = (f155 >= `INH(p150)) ? `INH(p150) : f155;
        f155 = (f155 >= `INH(p152)) ? `INH(p152) : f155;
        f155 = (f155 > p153) ? p153 : f155;
        f156 = 131071;
        f156 = (f156 > p16) ? p16 : f156;
        f156 = (f156 >= `INH(p155)) ? `INH(p155) : f156;
        f157 = 131071;
        f157 = (f157 > p154) ? p154 : f157;
        f157 = (f157 >= `INH(p156)) ? `INH(p156) : f157;
        f158 = 131071;
        f158 = (f158 >= `INH(p16)) ? `INH(p16) : f158;
        f158 = (f158 >= `INH(p155)) ? `INH(p155) : f158;
        f158 = (f158 > p156) ? p156 : f158;
        f159 = 131071;
        f159 = (f159 >= `INH(p154)) ? `INH(p154) : f159;
        f159 = (f159 >= `INH(p156)) ? `INH(p156) : f159;
        f159 = (f159 > p157) ? p157 : f159;
        f160 = 131071;
        f160 = (f160 > p21) ? p21 : f160;
        f160 = (f160 >= `INH(p159)) ? `INH(p159) : f160;
        f161 = 131071;
        f161 = (f161 > p158) ? p158 : f161;
        f161 = (f161 >= `INH(p160)) ? `INH(p160) : f161;
        f162 = 131071;
        f162 = (f162 >= `INH(p21)) ? `INH(p21) : f162;
        f162 = (f162 >= `INH(p159)) ? `INH(p159) : f162;
        f162 = (f162 > p160) ? p160 : f162;
        f163 = 131071;
        f163 = (f163 >= `INH(p158)) ? `INH(p158) : f163;
        f163 = (f163 >= `INH(p160)) ? `INH(p160) : f163;
        f163 = (f163 > p161) ? p161 : f163;
        f164 = 131071;
        f164 = (f164 >= `INH(p5)) ? `INH(p5) : f164;
        f164 = (f164 > p155) ? p155 : f164;
        f164 = (f164 > p159) ? p159 : f164;
        f165 = 131071;
        f165 = (f165 > p152) ? p152 : f165;
        f165 = (f165 >= `INH(p157)) ? `INH(p157) : f165;
        f165 = (f165 >= `INH(p161)) ? `INH(p161) : f165;
        f166 = 131071;
        f166 = (f166 > p151) ? p151 : f166;
        f166 = (f166 >= `INH(p162)) ? `INH(p162) : f166;
        f167 = 131071;
        f167 = (f167 > p22) ? p22 : f167;
        f167 = (f167 >= `INH(p153)) ? `INH(p153) : f167;
        f168 = 131071;
        f168 = (f168 >= `INH(p22)) ? `INH(p22) : f168;
        f168 = (f168 >= `INH(p153)) ? `INH(p153) : f168;
        f168 = (f168 > p162) ? p162 : f168;
        f169 = 131071;
        f169 = (f169 > p6) ? p6 : f169;
        f169 = (f169 >= `INH(p151)) ? `INH(p151) : f169;
        f169 = (f169 >= `INH(p162)) ? `INH(p162) : f169;
        f170 = 131071;
        f170 = (f170 >= `INH(p164)) ? `INH(p164) : f170;
        f170 = (f170 >= `INH(p165)) ? `INH(p165) : f170;
        f170 = (f170 > p169) ? p169 : f170;
        f171 = 131071;
        f171 = (f171 > p163) ? p163 : f171;
        f171 = (f171 >= `INH(p169)) ? `INH(p169) : f171;
        f172 = 131071;
        f172 = (f172 > p167) ? p167 : f172;
        f172 = (f172 >= `INH(p169)) ? `INH(p169) : f172;
        f173 = 131071;
        f173 = (f173 >= p164/2) ? p164/2 : f173;
        f173 = (f173 >= `INH(p168)) ? `INH(p168) : f173;
        f174 = 131071;
        f174 = (f174 >= `INH(p168)) ? `INH(p168) : f174;
        f174 = (f174 > p171) ? p171 : f174;
        f175 = 131071;
        f175 = (f175 > p164) ? p164 : f175;
        f175 = (f175 >= `INH(p171)) ? `INH(p171) : f175;
        f175 = (f175 > p173) ? p173 : f175;
        f176 = 131071;
        f176 = (f176 >= `INH(p171)) ? `INH(p171) : f176;
        f176 = (f176 > p174) ? p174 : f176;
        f177 = 131071;
        f177 = (f177 > p163) ? p163 : f177;
        f177 = (f177 >= `INH(p173)) ? `INH(p173) : f177;
        f177 = (f177 >= `INH(p174)) ? `INH(p174) : f177;
        f178 = 131071;
        f178 = (f178 > p163) ? p163 : f178;
        f178 = (f178 >= `INH(p172)) ? `INH(p172) : f178;
        f178 = (f178 >= `INH(p174)) ? `INH(p174) : f178;
        f179 = 131071;
        f179 = (f179 >= `INH(p174)) ? `INH(p174) : f179;
        f179 = (f179 > p176) ? p176 : f179;
        f180 = 131071;
        f180 = (f180 > p170) ? p170 : f180;
        f180 = (f180 >= `INH(p176)) ? `INH(p176) : f180;
        f181 = 131071;
        f181 = (f181 >= `INH(p176)) ? `INH(p176) : f181;
        f181 = (f181 > p177) ? p177 : f181;
        f182 = 131071;
        f182 = (f182 > p175) ? p175 : f182;
        f182 = (f182 >= `INH(p177)) ? `INH(p177) : f182;
        f183 = 131071;
        f183 = (f183 > p165) ? p165 : f183;
        f183 = (f183 > p172) ? p172 : f183;
        f183 = (f183 >= `INH(p173)) ? `INH(p173) : f183;
        f183 = (f183 >= `INH(p177)) ? `INH(p177) : f183;
        f184 = 131071;
        f184 = (f184 > p165) ? p165 : f184;
        f184 = (f184 >= `INH(p172)) ? `INH(p172) : f184;
        f184 = (f184 >= `INH(p177)) ? `INH(p177) : f184;
        f185 = 131071;
        f185 = (f185 > p23) ? p23 : f185;
        f185 = (f185 >= `INH(p179)) ? `INH(p179) : f185;
        f186 = 131071;
        f186 = (f186 > p178) ? p178 : f186;
        f186 = (f186 >= `INH(p180)) ? `INH(p180) : f186;
        f187 = 131071;
        f187 = (f187 >= `INH(p23)) ? `INH(p23) : f187;
        f187 = (f187 >= `INH(p179)) ? `INH(p179) : f187;
        f187 = (f187 > p180) ? p180 : f187;
        f188 = 131071;
        f188 = (f188 >= `INH(p178)) ? `INH(p178) : f188;
        f188 = (f188 >= `INH(p180)) ? `INH(p180) : f188;
        f188 = (f188 > p181) ? p181 : f188;
        f189 = 131071;
        f189 = (f189 > p24) ? p24 : f189;
        f189 = (f189 >= `INH(p183)) ? `INH(p183) : f189;
        f190 = 131071;
        f190 = (f190 > p182) ? p182 : f190;
        f190 = (f190 >= `INH(p184)) ? `INH(p184) : f190;
        f191 = 131071;
        f191 = (f191 >= `INH(p24)) ? `INH(p24) : f191;
        f191 = (f191 >= `INH(p183)) ? `INH(p183) : f191;
        f191 = (f191 > p184) ? p184 : f191;
        f192 = 131071;
        f192 = (f192 >= `INH(p182)) ? `INH(p182) : f192;
        f192 = (f192 >= `INH(p184)) ? `INH(p184) : f192;
        f192 = (f192 > p185) ? p185 : f192;
        f193 = 131071;
        f193 = (f193 >= `INH(p6)) ? `INH(p6) : f193;
        f193 = (f193 > p179) ? p179 : f193;
        f193 = (f193 > p183) ? p183 : f193;
        f194 = 131071;
        f194 = (f194 > p165) ? p165 : f194;
        f194 = (f194 >= `INH(p181)) ? `INH(p181) : f194;
        f194 = (f194 >= `INH(p185)) ? `INH(p185) : f194;
        f195 = 131071;
        f195 = (f195 > p166) ? p166 : f195;
        f195 = (f195 >= `INH(p186)) ? `INH(p186) : f195;
        f196 = 131071;
        f196 = (f196 > p25) ? p25 : f196;
        f196 = (f196 >= `INH(p167)) ? `INH(p167) : f196;
        f197 = 131071;
        f197 = (f197 >= `INH(p25)) ? `INH(p25) : f197;
        f197 = (f197 >= `INH(p167)) ? `INH(p167) : f197;
        f197 = (f197 > p186) ? p186 : f197;
        f198 = 131071;
        f198 = (f198 > p7) ? p7 : f198;
        f198 = (f198 >= `INH(p166)) ? `INH(p166) : f198;
        f198 = (f198 >= `INH(p186)) ? `INH(p186) : f198;
        f199 = 131071;
        f199 = (f199 > p188) ? p188 : f199;
        f199 = (f199 >= `INH(p190)) ? `INH(p190) : f199;
        f200 = 131071;
        f200 = (f200 >= `INH(p187)) ? `INH(p187) : f200;
        f200 = (f200 >= `INH(p188)) ? `INH(p188) : f200;
        f200 = (f200 >= `INH(p190)) ? `INH(p190) : f200;
        f200 = (f200 > p191) ? p191 : f200;
        f201 = 131071;
        f201 = (f201 > p25) ? p25 : f201;
        f201 = (f201 >= `INH(p193)) ? `INH(p193) : f201;
        f202 = 131071;
        f202 = (f202 > p192) ? p192 : f202;
        f202 = (f202 >= `INH(p194)) ? `INH(p194) : f202;
        f203 = 131071;
        f203 = (f203 >= `INH(p25)) ? `INH(p25) : f203;
        f203 = (f203 >= `INH(p193)) ? `INH(p193) : f203;
        f203 = (f203 > p194) ? p194 : f203;
        f204 = 131071;
        f204 = (f204 >= `INH(p192)) ? `INH(p192) : f204;
        f204 = (f204 >= `INH(p194)) ? `INH(p194) : f204;
        f204 = (f204 > p195) ? p195 : f204;
        f205 = 131071;
        f205 = (f205 > p22) ? p22 : f205;
        f205 = (f205 >= `INH(p197)) ? `INH(p197) : f205;
        f206 = 131071;
        f206 = (f206 > p196) ? p196 : f206;
        f206 = (f206 >= `INH(p198)) ? `INH(p198) : f206;
        f207 = 131071;
        f207 = (f207 >= `INH(p22)) ? `INH(p22) : f207;
        f207 = (f207 >= `INH(p197)) ? `INH(p197) : f207;
        f207 = (f207 > p198) ? p198 : f207;
        f208 = 131071;
        f208 = (f208 >= `INH(p196)) ? `INH(p196) : f208;
        f208 = (f208 >= `INH(p198)) ? `INH(p198) : f208;
        f208 = (f208 > p199) ? p199 : f208;
        f209 = 131071;
        f209 = (f209 >= `INH(p7)) ? `INH(p7) : f209;
        f209 = (f209 > p193) ? p193 : f209;
        f209 = (f209 > p197) ? p197 : f209;
        f210 = 131071;
        f210 = (f210 > p190) ? p190 : f210;
        f210 = (f210 >= `INH(p195)) ? `INH(p195) : f210;
        f210 = (f210 >= `INH(p199)) ? `INH(p199) : f210;
        f211 = 131071;
        f211 = (f211 > p189) ? p189 : f211;
        f211 = (f211 >= `INH(p200)) ? `INH(p200) : f211;
        f212 = 131071;
        f212 = (f212 > p26) ? p26 : f212;
        f212 = (f212 >= `INH(p191)) ? `INH(p191) : f212;
        f213 = 131071;
        f213 = (f213 >= `INH(p26)) ? `INH(p26) : f213;
        f213 = (f213 >= `INH(p191)) ? `INH(p191) : f213;
        f213 = (f213 > p200) ? p200 : f213;
        f214 = 131071;
        f214 = (f214 > p8) ? p8 : f214;
        f214 = (f214 >= `INH(p189)) ? `INH(p189) : f214;
        f214 = (f214 >= `INH(p200)) ? `INH(p200) : f214;
        f215 = 131071;
        f215 = (f215 > p202) ? p202 : f215;
        f215 = (f215 >= `INH(p204)) ? `INH(p204) : f215;
        f216 = 131071;
        f216 = (f216 >= `INH(p201)) ? `INH(p201) : f216;
        f216 = (f216 >= `INH(p202)) ? `INH(p202) : f216;
        f216 = (f216 >= `INH(p204)) ? `INH(p204) : f216;
        f216 = (f216 > p205) ? p205 : f216;
        f217 = 131071;
        f217 = (f217 > p26) ? p26 : f217;
        f217 = (f217 >= `INH(p207)) ? `INH(p207) : f217;
        f218 = 131071;
        f218 = (f218 > p206) ? p206 : f218;
        f218 = (f218 >= `INH(p208)) ? `INH(p208) : f218;
        f219 = 131071;
        f219 = (f219 >= `INH(p26)) ? `INH(p26) : f219;
        f219 = (f219 >= `INH(p207)) ? `INH(p207) : f219;
        f219 = (f219 > p208) ? p208 : f219;
        f220 = 131071;
        f220 = (f220 >= `INH(p206)) ? `INH(p206) : f220;
        f220 = (f220 >= `INH(p208)) ? `INH(p208) : f220;
        f220 = (f220 > p209) ? p209 : f220;
        f221 = 131071;
        f221 = (f221 > p27) ? p27 : f221;
        f221 = (f221 >= `INH(p211)) ? `INH(p211) : f221;
        f222 = 131071;
        f222 = (f222 > p210) ? p210 : f222;
        f222 = (f222 >= `INH(p212)) ? `INH(p212) : f222;
        f223 = 131071;
        f223 = (f223 >= `INH(p27)) ? `INH(p27) : f223;
        f223 = (f223 >= `INH(p211)) ? `INH(p211) : f223;
        f223 = (f223 > p212) ? p212 : f223;
        f224 = 131071;
        f224 = (f224 >= `INH(p210)) ? `INH(p210) : f224;
        f224 = (f224 >= `INH(p212)) ? `INH(p212) : f224;
        f224 = (f224 > p213) ? p213 : f224;
        f225 = 131071;
        f225 = (f225 >= `INH(p8)) ? `INH(p8) : f225;
        f225 = (f225 > p207) ? p207 : f225;
        f225 = (f225 > p211) ? p211 : f225;
        f226 = 131071;
        f226 = (f226 > p204) ? p204 : f226;
        f226 = (f226 >= `INH(p209)) ? `INH(p209) : f226;
        f226 = (f226 >= `INH(p213)) ? `INH(p213) : f226;
        f227 = 131071;
        f227 = (f227 > p203) ? p203 : f227;
        f227 = (f227 >= `INH(p214)) ? `INH(p214) : f227;
        f228 = 131071;
        f228 = (f228 > p28) ? p28 : f228;
        f228 = (f228 >= `INH(p205)) ? `INH(p205) : f228;
        f229 = 131071;
        f229 = (f229 >= `INH(p28)) ? `INH(p28) : f229;
        f229 = (f229 >= `INH(p205)) ? `INH(p205) : f229;
        f229 = (f229 > p214) ? p214 : f229;
        f230 = 131071;
        f230 = (f230 > p9) ? p9 : f230;
        f230 = (f230 >= `INH(p203)) ? `INH(p203) : f230;
        f230 = (f230 >= `INH(p214)) ? `INH(p214) : f230;
        if(f9>0)
                f0 = 0;
        if(f10>0)
                f11 = 0;
        if(f12>0)
                f13 = 0;
        if(f14>0)
                f15 = 0;
        if(f16>0)
                f18 = 0;
        if(f17>0)
                f18 = 0;
        if(f19>0)
                f20 = 0;
        if(f21>0)
                f22 = 0;
        if(f21>0)
                f23 = 0;
        if(f38>0)
                f1 = 0;
        if(f39>0)
                f40 = 0;
        if(f41>0)
                f42 = 0;
        if(f43>0)
                f44 = 0;
        if(f45>0)
                f47 = 0;
        if(f46>0)
                f47 = 0;
        if(f48>0)
                f49 = 0;
        if(f50>0)
                f51 = 0;
        if(f50>0)
                f52 = 0;
        if(f67>0)
                f2 = 0;
        if(f68>0)
                f69 = 0;
        if(f70>0)
                f71 = 0;
        if(f72>0)
                f73 = 0;
        if(f74>0)
                f76 = 0;
        if(f75>0)
                f76 = 0;
        if(f77>0)
                f78 = 0;
        if(f79>0)
                f80 = 0;
        if(f79>0)
                f81 = 0;
        if(f96>0)
                f3 = 0;
        if(f97>0)
                f98 = 0;
        if(f99>0)
                f100 = 0;
        if(f101>0)
                f102 = 0;
        if(f103>0)
                f105 = 0;
        if(f104>0)
                f105 = 0;
        if(f106>0)
                f107 = 0;
        if(f108>0)
                f109 = 0;
        if(f108>0)
                f110 = 0;
        if(f125>0)
                f4 = 0;
        if(f126>0)
                f127 = 0;
        if(f128>0)
                f129 = 0;
        if(f130>0)
                f131 = 0;
        if(f132>0)
                f134 = 0;
        if(f133>0)
                f134 = 0;
        if(f135>0)
                f136 = 0;
        if(f137>0)
                f138 = 0;
        if(f137>0)
                f139 = 0;
        if(f170>0)
                f6 = 0;
        if(f171>0)
                f172 = 0;
        if(f173>0)
                f174 = 0;
        if(f175>0)
                f176 = 0;
        if(f177>0)
                f179 = 0;
        if(f178>0)
                f179 = 0;
        if(f180>0)
                f181 = 0;
        if(f182>0)
                f183 = 0;
        if(f182>0)
                f184 = 0;
        tf = (f0>0)?1:(f1>0)?2:(f2>0)?3:(f3>0)?4:(f4>0)?5:(f5>0)?6:(f6>0)?7:(f7>0)?8:(f8>0)?9:(f9>0)?10:(f10>0)?11:(f11>0)?12:(f12>0)?13:(f13>0)?14:(f14>0)?15:(f15>0)?16:(f16>0)?17:(f17>0)?18:(f18>0)?19:(f19>0)?20:(f20>0)?21:(f21>0)?22:(f22>0)?23:(f23>0)?24:(f24>0)?25:(f25>0)?26:(f26>0)?27:(f27>0)?28:(f28>0)?29:(f29>0)?30:(f30>0)?31:(f31>0)?32:(f32>0)?33:(f33>0)?34:(f34>0)?35:(f35>0)?36:(f36>0)?37:(f37>0)?38:(f38>0)?39:(f39>0)?40:(f40>0)?41:(f41>0)?42:(f42>0)?43:(f43>0)?44:(f44>0)?45:(f45>0)?46:(f46>0)?47:(f47>0)?48:(f48>0)?49:(f49>0)?50:(f50>0)?51:(f51>0)?52:(f52>0)?53:(f53>0)?54:(f54>0)?55:(f55>0)?56:(f56>0)?57:(f57>0)?58:(f58>0)?59:(f59>0)?60:(f60>0)?61:(f61>0)?62:(f62>0)?63:(f63>0)?64:(f64>0)?65:(f65>0)?66:(f66>0)?67:(f67>0)?68:(f68>0)?69:(f69>0)?70:(f70>0)?71:(f71>0)?72:(f72>0)?73:(f73>0)?74:(f74>0)?75:(f75>0)?76:(f76>0)?77:(f77>0)?78:(f78>0)?79:(f79>0)?80:(f80>0)?81:(f81>0)?82:(f82>0)?83:(f83>0)?84:(f84>0)?85:(f85>0)?86:(f86>0)?87:(f87>0)?88:(f88>0)?89:(f89>0)?90:(f90>0)?91:(f91>0)?92:(f92>0)?93:(f93>0)?94:(f94>0)?95:(f95>0)?96:(f96>0)?97:(f97>0)?98:(f98>0)?99:(f99>0)?100:(f100>0)?101:(f101>0)?102:(f102>0)?103:(f103>0)?104:(f104>0)?105:(f105>0)?106:(f106>0)?107:(f107>0)?108:(f108>0)?109:(f109>0)?110:(f110>0)?111:(f111>0)?112:(f112>0)?113:(f113>0)?114:(f114>0)?115:(f115>0)?116:(f116>0)?117:(f117>0)?118:(f118>0)?119:(f119>0)?120:(f120>0)?121:(f121>0)?122:(f122>0)?123:(f123>0)?124:(f124>0)?125:(f125>0)?126:(f126>0)?127:(f127>0)?128:(f128>0)?129:(f129>0)?130:(f130>0)?131:(f131>0)?132:(f132>0)?133:(f133>0)?134:(f134>0)?135:(f135>0)?136:(f136>0)?137:(f137>0)?138:(f138>0)?139:(f139>0)?140:(f140>0)?141:(f141>0)?142:(f142>0)?143:(f143>0)?144:(f144>0)?145:(f145>0)?146:(f146>0)?147:(f147>0)?148:(f148>0)?149:(f149>0)?150:(f150>0)?151:(f151>0)?152:(f152>0)?153:(f153>0)?154:(f154>0)?155:(f155>0)?156:(f156>0)?157:(f157>0)?158:(f158>0)?159:(f159>0)?160:(f160>0)?161:(f161>0)?162:(f162>0)?163:(f163>0)?164:(f164>0)?165:(f165>0)?166:(f166>0)?167:(f167>0)?168:(f168>0)?169:(f169>0)?170:(f170>0)?171:(f171>0)?172:(f172>0)?173:(f173>0)?174:(f174>0)?175:(f175>0)?176:(f176>0)?177:(f177>0)?178:(f178>0)?179:(f179>0)?180:(f180>0)?181:(f181>0)?182:(f182>0)?183:(f183>0)?184:(f184>0)?185:(f185>0)?186:(f186>0)?187:(f187>0)?188:(f188>0)?189:(f189>0)?190:(f190>0)?191:(f191>0)?192:(f192>0)?193:(f193>0)?194:(f194>0)?195:(f195>0)?196:(f196>0)?197:(f197>0)?198:(f198>0)?199:(f199>0)?200:(f200>0)?201:(f201>0)?202:(f202>0)?203:(f203>0)?204:(f204>0)?205:(f205>0)?206:(f206>0)?207:(f207>0)?208:(f208>0)?209:(f209>0)?210:(f210>0)?211:(f211>0)?212:(f212>0)?213:(f213>0)?214:(f214>0)?215:(f215>0)?216:(f216>0)?217:(f217>0)?218:(f218>0)?219:(f219>0)?220:(f220>0)?221:(f221>0)?222:(f222>0)?223:(f223>0)?224:(f224>0)?225:(f225>0)?226:(f226>0)?227:(f227>0)?228:(f228>0)?229:(f229>0)?230:(f230>0)?231:0;
        case(tf)
                1: begin
                        tc = f0;
                        p34 = p34 - tc;
                        p31 = p31 + tc;
                end
                2: begin
                        tc = f1;
                        p58 = p58 - tc;
                        p55 = p55 + tc;
                end
                3: begin
                        tc = f2;
                        p82 = p82 - tc;
                        p79 = p79 + tc;
                end
                4: begin
                        tc = f3;
                        p106 = p106 - tc;
                        p103 = p103 + tc;
                end
                5: begin
                        tc = f4;
                        p130 = p130 - tc;
                        p127 = p127 + tc;
                end
                6: begin
                        tc = f5;
                        p149 = p149 - tc;
                        p151 = p151 + tc;
                end
                7: begin
                        tc = f6;
                        p168 = p168 - tc;
                        p165 = p165 + tc;
                end
                8: begin
                        tc = f7;
                        p187 = p187 - tc;
                        p189 = p189 + tc;
                end
                9: begin
                        tc = f8;
                        p201 = p201 - tc;
                        p203 = p203 + tc;
                end
                10: begin
                        tc = f9;
                        p35 = p35 - tc;
                        p31 = p31 + tc;
                end
                11: begin
                        tc = f10;
                        p29 = p29 - tc;
                end
                12: begin
                        tc = f11;
                        p33 = p33 - tc;
                        p35 = p35 + tc;
                end
                13: begin
                        tc = f12;
                        p30 = p30 - tc*2;
                        p36 = p36 + tc;
                end
                14: begin
                        tc = f13;
                        p37 = p37 - tc;
                        p34 = p34 + tc;
                end
                15: begin
                        tc = f14;
                        p30 = p30 - tc;
                        p39 = p39 - tc;
                        p38 = p38 + tc;
                end
                16: begin
                        tc = f15;
                        p40 = p40 - tc;
                        p37 = p37 + tc;
                end
                17: begin
                        tc = f16;
                        p29 = p29 - tc;
                        p32 = p32 + tc;
                        p41 = p41 + tc;
                end
                18: begin
                        tc = f17;
                        p29 = p29 - tc;
                        p41 = p41 + tc;
                end
                19: begin
                        tc = f18;
                        p42 = p42 - tc;
                        p40 = p40 + tc;
                end
                20: begin
                        tc = f19;
                        p36 = p36 - tc;
                        p30 = p30 + tc;
                end
                21: begin
                        tc = f20;
                        p43 = p43 - tc;
                        p42 = p42 + tc;
                end
                22: begin
                        tc = f21;
                        p41 = p41 - tc;
                        p29 = p29 + tc*2;
                end
                23: begin
                        tc = f22;
                        p31 = p31 - tc;
                        p38 = p38 - tc;
                        p39 = p39 + tc;
                        p43 = p43 + tc;
                end
                24: begin
                        tc = f23;
                        p31 = p31 - tc;
                        p43 = p43 + tc;
                end
                25: begin
                        tc = f24;
                        p10 = p10 - tc;
                        p29 = p29 + tc;
                        p44 = p44 + tc;
                end
                26: begin
                        tc = f25;
                        p44 = p44 - tc;
                        p10 = p10 + tc;
                end
                27: begin
                        tc = f26;
                        p46 = p46 - tc;
                        p45 = p45 + tc;
                end
                28: begin
                        tc = f27;
                        p47 = p47 - tc;
                        p46 = p46 + tc;
                end
                29: begin
                        tc = f28;
                        p11 = p11 - tc;
                        p30 = p30 + tc;
                        p48 = p48 + tc;
                end
                30: begin
                        tc = f29;
                        p48 = p48 - tc;
                        p11 = p11 + tc;
                end
                31: begin
                        tc = f30;
                        p50 = p50 - tc;
                        p49 = p49 + tc;
                end
                32: begin
                        tc = f31;
                        p51 = p51 - tc;
                        p50 = p50 + tc;
                end
                33: begin
                        tc = f32;
                        p45 = p45 - tc;
                        p49 = p49 - tc;
                        p0 = p0 + tc;
                end
                34: begin
                        tc = f33;
                        p31 = p31 - tc;
                        p47 = p47 + tc;
                        p51 = p51 + tc;
                end
                35: begin
                        tc = f34;
                        p32 = p32 - tc;
                        p12 = p12 + tc;
                end
                36: begin
                        tc = f35;
                        p12 = p12 - tc;
                end
                37: begin
                        tc = f36;
                        p52 = p52 - tc;
                        p33 = p33 + tc;
                end
                38: begin
                        tc = f37;
                        p1 = p1 - tc;
                        p52 = p52 + tc;
                end
                39: begin
                        tc = f38;
                        p59 = p59 - tc;
                        p55 = p55 + tc;
                end
                40: begin
                        tc = f39;
                        p53 = p53 - tc;
                end
                41: begin
                        tc = f40;
                        p57 = p57 - tc;
                        p59 = p59 + tc;
                end
                42: begin
                        tc = f41;
                        p54 = p54 - tc*2;
                        p60 = p60 + tc;
                end
                43: begin
                        tc = f42;
                        p61 = p61 - tc;
                        p58 = p58 + tc;
                end
                44: begin
                        tc = f43;
                        p54 = p54 - tc;
                        p63 = p63 - tc;
                        p62 = p62 + tc;
                end
                45: begin
                        tc = f44;
                        p64 = p64 - tc;
                        p61 = p61 + tc;
                end
                46: begin
                        tc = f45;
                        p53 = p53 - tc;
                        p56 = p56 + tc;
                        p65 = p65 + tc;
                end
                47: begin
                        tc = f46;
                        p53 = p53 - tc;
                        p65 = p65 + tc;
                end
                48: begin
                        tc = f47;
                        p66 = p66 - tc;
                        p64 = p64 + tc;
                end
                49: begin
                        tc = f48;
                        p60 = p60 - tc;
                        p54 = p54 + tc;
                end
                50: begin
                        tc = f49;
                        p67 = p67 - tc;
                        p66 = p66 + tc;
                end
                51: begin
                        tc = f50;
                        p65 = p65 - tc;
                        p53 = p53 + tc*2;
                end
                52: begin
                        tc = f51;
                        p55 = p55 - tc;
                        p62 = p62 - tc;
                        p63 = p63 + tc;
                        p67 = p67 + tc;
                end
                53: begin
                        tc = f52;
                        p55 = p55 - tc;
                        p67 = p67 + tc;
                end
                54: begin
                        tc = f53;
                        p12 = p12 - tc;
                        p53 = p53 + tc;
                        p68 = p68 + tc;
                end
                55: begin
                        tc = f54;
                        p68 = p68 - tc;
                        p12 = p12 + tc;
                end
                56: begin
                        tc = f55;
                        p70 = p70 - tc;
                        p69 = p69 + tc;
                end
                57: begin
                        tc = f56;
                        p71 = p71 - tc;
                        p70 = p70 + tc;
                end
                58: begin
                        tc = f57;
                        p13 = p13 - tc;
                        p54 = p54 + tc;
                        p72 = p72 + tc;
                end
                59: begin
                        tc = f58;
                        p72 = p72 - tc;
                        p13 = p13 + tc;
                end
                60: begin
                        tc = f59;
                        p74 = p74 - tc;
                        p73 = p73 + tc;
                end
                61: begin
                        tc = f60;
                        p75 = p75 - tc;
                        p74 = p74 + tc;
                end
                62: begin
                        tc = f61;
                        p69 = p69 - tc;
                        p73 = p73 - tc;
                        p1 = p1 + tc;
                end
                63: begin
                        tc = f62;
                        p55 = p55 - tc;
                        p71 = p71 + tc;
                        p75 = p75 + tc;
                end
                64: begin
                        tc = f63;
                        p56 = p56 - tc;
                        p14 = p14 + tc;
                end
                65: begin
                        tc = f64;
                        p14 = p14 - tc;
                end
                66: begin
                        tc = f65;
                        p76 = p76 - tc;
                        p57 = p57 + tc;
                end
                67: begin
                        tc = f66;
                        p2 = p2 - tc;
                        p76 = p76 + tc;
                end
                68: begin
                        tc = f67;
                        p83 = p83 - tc;
                        p79 = p79 + tc;
                end
                69: begin
                        tc = f68;
                        p77 = p77 - tc;
                end
                70: begin
                        tc = f69;
                        p81 = p81 - tc;
                        p83 = p83 + tc;
                end
                71: begin
                        tc = f70;
                        p78 = p78 - tc*2;
                        p84 = p84 + tc;
                end
                72: begin
                        tc = f71;
                        p85 = p85 - tc;
                        p82 = p82 + tc;
                end
                73: begin
                        tc = f72;
                        p78 = p78 - tc;
                        p87 = p87 - tc;
                        p86 = p86 + tc;
                end
                74: begin
                        tc = f73;
                        p88 = p88 - tc;
                        p85 = p85 + tc;
                end
                75: begin
                        tc = f74;
                        p77 = p77 - tc;
                        p80 = p80 + tc;
                        p89 = p89 + tc;
                end
                76: begin
                        tc = f75;
                        p77 = p77 - tc;
                        p89 = p89 + tc;
                end
                77: begin
                        tc = f76;
                        p90 = p90 - tc;
                        p88 = p88 + tc;
                end
                78: begin
                        tc = f77;
                        p84 = p84 - tc;
                        p78 = p78 + tc;
                end
                79: begin
                        tc = f78;
                        p91 = p91 - tc;
                        p90 = p90 + tc;
                end
                80: begin
                        tc = f79;
                        p89 = p89 - tc;
                        p77 = p77 + tc*2;
                end
                81: begin
                        tc = f80;
                        p79 = p79 - tc;
                        p86 = p86 - tc;
                        p87 = p87 + tc;
                        p91 = p91 + tc;
                end
                82: begin
                        tc = f81;
                        p79 = p79 - tc;
                        p91 = p91 + tc;
                end
                83: begin
                        tc = f82;
                        p14 = p14 - tc;
                        p77 = p77 + tc;
                        p92 = p92 + tc;
                end
                84: begin
                        tc = f83;
                        p92 = p92 - tc;
                        p14 = p14 + tc;
                end
                85: begin
                        tc = f84;
                        p94 = p94 - tc;
                        p93 = p93 + tc;
                end
                86: begin
                        tc = f85;
                        p95 = p95 - tc;
                        p94 = p94 + tc;
                end
                87: begin
                        tc = f86;
                        p15 = p15 - tc;
                        p78 = p78 + tc;
                        p96 = p96 + tc;
                end
                88: begin
                        tc = f87;
                        p96 = p96 - tc;
                        p15 = p15 + tc;
                end
                89: begin
                        tc = f88;
                        p98 = p98 - tc;
                        p97 = p97 + tc;
                end
                90: begin
                        tc = f89;
                        p99 = p99 - tc;
                        p98 = p98 + tc;
                end
                91: begin
                        tc = f90;
                        p93 = p93 - tc;
                        p97 = p97 - tc;
                        p2 = p2 + tc;
                end
                92: begin
                        tc = f91;
                        p79 = p79 - tc;
                        p95 = p95 + tc;
                        p99 = p99 + tc;
                end
                93: begin
                        tc = f92;
                        p80 = p80 - tc;
                        p16 = p16 + tc;
                end
                94: begin
                        tc = f93;
                        p16 = p16 - tc;
                end
                95: begin
                        tc = f94;
                        p100 = p100 - tc;
                        p81 = p81 + tc;
                end
                96: begin
                        tc = f95;
                        p3 = p3 - tc;
                        p100 = p100 + tc;
                end
                97: begin
                        tc = f96;
                        p107 = p107 - tc;
                        p103 = p103 + tc;
                end
                98: begin
                        tc = f97;
                        p101 = p101 - tc;
                end
                99: begin
                        tc = f98;
                        p105 = p105 - tc;
                        p107 = p107 + tc;
                end
                100: begin
                        tc = f99;
                        p102 = p102 - tc*2;
                        p108 = p108 + tc;
                end
                101: begin
                        tc = f100;
                        p109 = p109 - tc;
                        p106 = p106 + tc;
                end
                102: begin
                        tc = f101;
                        p102 = p102 - tc;
                        p111 = p111 - tc;
                        p110 = p110 + tc;
                end
                103: begin
                        tc = f102;
                        p112 = p112 - tc;
                        p109 = p109 + tc;
                end
                104: begin
                        tc = f103;
                        p101 = p101 - tc;
                        p104 = p104 + tc;
                        p113 = p113 + tc;
                end
                105: begin
                        tc = f104;
                        p101 = p101 - tc;
                        p113 = p113 + tc;
                end
                106: begin
                        tc = f105;
                        p114 = p114 - tc;
                        p112 = p112 + tc;
                end
                107: begin
                        tc = f106;
                        p108 = p108 - tc;
                        p102 = p102 + tc;
                end
                108: begin
                        tc = f107;
                        p115 = p115 - tc;
                        p114 = p114 + tc;
                end
                109: begin
                        tc = f108;
                        p113 = p113 - tc;
                        p101 = p101 + tc*2;
                end
                110: begin
                        tc = f109;
                        p103 = p103 - tc;
                        p110 = p110 - tc;
                        p111 = p111 + tc;
                        p115 = p115 + tc;
                end
                111: begin
                        tc = f110;
                        p103 = p103 - tc;
                        p115 = p115 + tc;
                end
                112: begin
                        tc = f111;
                        p17 = p17 - tc;
                        p101 = p101 + tc;
                        p116 = p116 + tc;
                end
                113: begin
                        tc = f112;
                        p116 = p116 - tc;
                        p17 = p17 + tc;
                end
                114: begin
                        tc = f113;
                        p118 = p118 - tc;
                        p117 = p117 + tc;
                end
                115: begin
                        tc = f114;
                        p119 = p119 - tc;
                        p118 = p118 + tc;
                end
                116: begin
                        tc = f115;
                        p18 = p18 - tc;
                        p102 = p102 + tc;
                        p120 = p120 + tc;
                end
                117: begin
                        tc = f116;
                        p120 = p120 - tc;
                        p18 = p18 + tc;
                end
                118: begin
                        tc = f117;
                        p122 = p122 - tc;
                        p121 = p121 + tc;
                end
                119: begin
                        tc = f118;
                        p123 = p123 - tc;
                        p122 = p122 + tc;
                end
                120: begin
                        tc = f119;
                        p117 = p117 - tc;
                        p121 = p121 - tc;
                        p3 = p3 + tc;
                end
                121: begin
                        tc = f120;
                        p103 = p103 - tc;
                        p119 = p119 + tc;
                        p123 = p123 + tc;
                end
                122: begin
                        tc = f121;
                        p104 = p104 - tc;
                        p19 = p19 + tc;
                end
                123: begin
                        tc = f122;
                        p19 = p19 - tc;
                end
                124: begin
                        tc = f123;
                        p124 = p124 - tc;
                        p105 = p105 + tc;
                end
                125: begin
                        tc = f124;
                        p4 = p4 - tc;
                        p124 = p124 + tc;
                end
                126: begin
                        tc = f125;
                        p131 = p131 - tc;
                        p127 = p127 + tc;
                end
                127: begin
                        tc = f126;
                        p125 = p125 - tc;
                end
                128: begin
                        tc = f127;
                        p129 = p129 - tc;
                        p131 = p131 + tc;
                end
                129: begin
                        tc = f128;
                        p126 = p126 - tc*2;
                        p132 = p132 + tc;
                end
                130: begin
                        tc = f129;
                        p133 = p133 - tc;
                        p130 = p130 + tc;
                end
                131: begin
                        tc = f130;
                        p126 = p126 - tc;
                        p135 = p135 - tc;
                        p134 = p134 + tc;
                end
                132: begin
                        tc = f131;
                        p136 = p136 - tc;
                        p133 = p133 + tc;
                end
                133: begin
                        tc = f132;
                        p125 = p125 - tc;
                        p128 = p128 + tc;
                        p137 = p137 + tc;
                end
                134: begin
                        tc = f133;
                        p125 = p125 - tc;
                        p137 = p137 + tc;
                end
                135: begin
                        tc = f134;
                        p138 = p138 - tc;
                        p136 = p136 + tc;
                end
                136: begin
                        tc = f135;
                        p132 = p132 - tc;
                        p126 = p126 + tc;
                end
                137: begin
                        tc = f136;
                        p139 = p139 - tc;
                        p138 = p138 + tc;
                end
                138: begin
                        tc = f137;
                        p137 = p137 - tc;
                        p125 = p125 + tc*2;
                end
                139: begin
                        tc = f138;
                        p127 = p127 - tc;
                        p134 = p134 - tc;
                        p135 = p135 + tc;
                        p139 = p139 + tc;
                end
                140: begin
                        tc = f139;
                        p127 = p127 - tc;
                        p139 = p139 + tc;
                end
                141: begin
                        tc = f140;
                        p19 = p19 - tc;
                        p125 = p125 + tc;
                        p140 = p140 + tc;
                end
                142: begin
                        tc = f141;
                        p140 = p140 - tc;
                        p19 = p19 + tc;
                end
                143: begin
                        tc = f142;
                        p142 = p142 - tc;
                        p141 = p141 + tc;
                end
                144: begin
                        tc = f143;
                        p143 = p143 - tc;
                        p142 = p142 + tc;
                end
                145: begin
                        tc = f144;
                        p20 = p20 - tc;
                        p126 = p126 + tc;
                        p144 = p144 + tc;
                end
                146: begin
                        tc = f145;
                        p144 = p144 - tc;
                        p20 = p20 + tc;
                end
                147: begin
                        tc = f146;
                        p146 = p146 - tc;
                        p145 = p145 + tc;
                end
                148: begin
                        tc = f147;
                        p147 = p147 - tc;
                        p146 = p146 + tc;
                end
                149: begin
                        tc = f148;
                        p141 = p141 - tc;
                        p145 = p145 - tc;
                        p4 = p4 + tc;
                end
                150: begin
                        tc = f149;
                        p127 = p127 - tc;
                        p143 = p143 + tc;
                        p147 = p147 + tc;
                end
                151: begin
                        tc = f150;
                        p128 = p128 - tc;
                        p21 = p21 + tc;
                end
                152: begin
                        tc = f151;
                        p21 = p21 - tc;
                end
                153: begin
                        tc = f152;
                        p148 = p148 - tc;
                        p129 = p129 + tc;
                end
                154: begin
                        tc = f153;
                        p5 = p5 - tc;
                        p148 = p148 + tc;
                end
                155: begin
                        tc = f154;
                        p150 = p150 - tc;
                        p151 = p151 + tc;
                end
                156: begin
                        tc = f155;
                        p153 = p153 - tc;
                        p152 = p152 + tc;
                end
                157: begin
                        tc = f156;
                        p16 = p16 - tc;
                        p149 = p149 + tc;
                        p154 = p154 + tc;
                end
                158: begin
                        tc = f157;
                        p154 = p154 - tc;
                        p16 = p16 + tc;
                end
                159: begin
                        tc = f158;
                        p156 = p156 - tc;
                        p155 = p155 + tc;
                end
                160: begin
                        tc = f159;
                        p157 = p157 - tc;
                        p156 = p156 + tc;
                end
                161: begin
                        tc = f160;
                        p21 = p21 - tc;
                        p150 = p150 + tc;
                        p158 = p158 + tc;
                end
                162: begin
                        tc = f161;
                        p158 = p158 - tc;
                        p21 = p21 + tc;
                end
                163: begin
                        tc = f162;
                        p160 = p160 - tc;
                        p159 = p159 + tc;
                end
                164: begin
                        tc = f163;
                        p161 = p161 - tc;
                        p160 = p160 + tc;
                end
                165: begin
                        tc = f164;
                        p155 = p155 - tc;
                        p159 = p159 - tc;
                        p5 = p5 + tc;
                end
                166: begin
                        tc = f165;
                        p152 = p152 - tc;
                        p157 = p157 + tc;
                        p161 = p161 + tc;
                end
                167: begin
                        tc = f166;
                        p151 = p151 - tc;
                        p22 = p22 + tc;
                end
                168: begin
                        tc = f167;
                        p22 = p22 - tc;
                end
                169: begin
                        tc = f168;
                        p162 = p162 - tc;
                        p153 = p153 + tc;
                end
                170: begin
                        tc = f169;
                        p6 = p6 - tc;
                        p162 = p162 + tc;
                end
                171: begin
                        tc = f170;
                        p169 = p169 - tc;
                        p165 = p165 + tc;
                end
                172: begin
                        tc = f171;
                        p163 = p163 - tc;
                end
                173: begin
                        tc = f172;
                        p167 = p167 - tc;
                        p169 = p169 + tc;
                end
                174: begin
                        tc = f173;
                        p164 = p164 - tc*2;
                        p170 = p170 + tc;
                end
                175: begin
                        tc = f174;
                        p171 = p171 - tc;
                        p168 = p168 + tc;
                end
                176: begin
                        tc = f175;
                        p164 = p164 - tc;
                        p173 = p173 - tc;
                        p172 = p172 + tc;
                end
                177: begin
                        tc = f176;
                        p174 = p174 - tc;
                        p171 = p171 + tc;
                end
                178: begin
                        tc = f177;
                        p163 = p163 - tc;
                        p166 = p166 + tc;
                        p175 = p175 + tc;
                end
                179: begin
                        tc = f178;
                        p163 = p163 - tc;
                        p175 = p175 + tc;
                end
                180: begin
                        tc = f179;
                        p176 = p176 - tc;
                        p174 = p174 + tc;
                end
                181: begin
                        tc = f180;
                        p170 = p170 - tc;
                        p164 = p164 + tc;
                end
                182: begin
                        tc = f181;
                        p177 = p177 - tc;
                        p176 = p176 + tc;
                end
                183: begin
                        tc = f182;
                        p175 = p175 - tc;
                        p163 = p163 + tc*2;
                end
                184: begin
                        tc = f183;
                        p165 = p165 - tc;
                        p172 = p172 - tc;
                        p173 = p173 + tc;
                        p177 = p177 + tc;
                end
                185: begin
                        tc = f184;
                        p165 = p165 - tc;
                        p177 = p177 + tc;
                end
                186: begin
                        tc = f185;
                        p23 = p23 - tc;
                        p163 = p163 + tc;
                        p178 = p178 + tc;
                end
                187: begin
                        tc = f186;
                        p178 = p178 - tc;
                        p23 = p23 + tc;
                end
                188: begin
                        tc = f187;
                        p180 = p180 - tc;
                        p179 = p179 + tc;
                end
                189: begin
                        tc = f188;
                        p181 = p181 - tc;
                        p180 = p180 + tc;
                end
                190: begin
                        tc = f189;
                        p24 = p24 - tc;
                        p164 = p164 + tc;
                        p182 = p182 + tc;
                end
                191: begin
                        tc = f190;
                        p182 = p182 - tc;
                        p24 = p24 + tc;
                end
                192: begin
                        tc = f191;
                        p184 = p184 - tc;
                        p183 = p183 + tc;
                end
                193: begin
                        tc = f192;
                        p185 = p185 - tc;
                        p184 = p184 + tc;
                end
                194: begin
                        tc = f193;
                        p179 = p179 - tc;
                        p183 = p183 - tc;
                        p6 = p6 + tc;
                end
                195: begin
                        tc = f194;
                        p165 = p165 - tc;
                        p181 = p181 + tc;
                        p185 = p185 + tc;
                end
                196: begin
                        tc = f195;
                        p166 = p166 - tc;
                        p25 = p25 + tc;
                end
                197: begin
                        tc = f196;
                        p25 = p25 - tc;
                end
                198: begin
                        tc = f197;
                        p186 = p186 - tc;
                        p167 = p167 + tc;
                end
                199: begin
                        tc = f198;
                        p7 = p7 - tc;
                        p186 = p186 + tc;
                end
                200: begin
                        tc = f199;
                        p188 = p188 - tc;
                        p189 = p189 + tc;
                end
                201: begin
                        tc = f200;
                        p191 = p191 - tc;
                        p190 = p190 + tc;
                end
                202: begin
                        tc = f201;
                        p25 = p25 - tc;
                        p187 = p187 + tc;
                        p192 = p192 + tc;
                end
                203: begin
                        tc = f202;
                        p192 = p192 - tc;
                        p25 = p25 + tc;
                end
                204: begin
                        tc = f203;
                        p194 = p194 - tc;
                        p193 = p193 + tc;
                end
                205: begin
                        tc = f204;
                        p195 = p195 - tc;
                        p194 = p194 + tc;
                end
                206: begin
                        tc = f205;
                        p22 = p22 - tc;
                        p188 = p188 + tc;
                        p196 = p196 + tc;
                end
                207: begin
                        tc = f206;
                        p196 = p196 - tc;
                        p22 = p22 + tc;
                end
                208: begin
                        tc = f207;
                        p198 = p198 - tc;
                        p197 = p197 + tc;
                end
                209: begin
                        tc = f208;
                        p199 = p199 - tc;
                        p198 = p198 + tc;
                end
                210: begin
                        tc = f209;
                        p193 = p193 - tc;
                        p197 = p197 - tc;
                        p7 = p7 + tc;
                end
                211: begin
                        tc = f210;
                        p190 = p190 - tc;
                        p195 = p195 + tc;
                        p199 = p199 + tc;
                end
                212: begin
                        tc = f211;
                        p189 = p189 - tc;
                        p26 = p26 + tc;
                end
                213: begin
                        tc = f212;
                        p26 = p26 - tc;
                end
                214: begin
                        tc = f213;
                        p200 = p200 - tc;
                        p191 = p191 + tc;
                end
                215: begin
                        tc = f214;
                        p8 = p8 - tc;
                        p200 = p200 + tc;
                end
                216: begin
                        tc = f215;
                        p202 = p202 - tc;
                        p203 = p203 + tc;
                end
                217: begin
                        tc = f216;
                        p205 = p205 - tc;
                        p204 = p204 + tc;
                end
                218: begin
                        tc = f217;
                        p26 = p26 - tc;
                        p201 = p201 + tc;
                        p206 = p206 + tc;
                end
                219: begin
                        tc = f218;
                        p206 = p206 - tc;
                        p26 = p26 + tc;
                end
                220: begin
                        tc = f219;
                        p208 = p208 - tc;
                        p207 = p207 + tc;
                end
                221: begin
                        tc = f220;
                        p209 = p209 - tc;
                        p208 = p208 + tc;
                end
                222: begin
                        tc = f221;
                        p27 = p27 - tc;
                        p202 = p202 + tc;
                        p210 = p210 + tc;
                end
                223: begin
                        tc = f222;
                        p210 = p210 - tc;
                        p27 = p27 + tc;
                end
                224: begin
                        tc = f223;
                        p212 = p212 - tc;
                        p211 = p211 + tc;
                end
                225: begin
                        tc = f224;
                        p213 = p213 - tc;
                        p212 = p212 + tc;
                end
                226: begin
                        tc = f225;
                        p207 = p207 - tc;
                        p211 = p211 - tc;
                        p8 = p8 + tc;
                end
                227: begin
                        tc = f226;
                        p204 = p204 - tc;
                        p209 = p209 + tc;
                        p213 = p213 + tc;
                end
                228: begin
                        tc = f227;
                        p203 = p203 - tc;
                        p28 = p28 + tc;
                end
                229: begin
                        tc = f228;
                        p28 = p28 - tc;
                end
                230: begin
                        tc = f229;
                        p214 = p214 - tc;
                        p205 = p205 + tc;
                end
                231: begin
                        tc = f230;
                        p9 = p9 - tc;
                        p214 = p214 + tc;
                end
                default:;
        endcase
//        led = ~p28[5:0];
  if(tf>0) counter1=counter1+1;
end
end
reg [32:0] counter;

always @(posedge clk) begin
    if (counter < 32'd2_7500_0000)       //delay
        counter <= counter + 1'b1;
    else
        counter <= 32'd0;
end

always @(posedge clk) begin
    if (counter == 32'd0)       
        led <= ~counter1[47:42];
    else if (counter == 32'd2500_0000)       
        led <= ~counter1[41:36];
    else if (counter == 32'd5000_0000)       
        led <= ~counter1[35:30];
    else if (counter == 32'd7500_0000)       
        led <= ~counter1[29:24];
    else if (counter == 32'd1_0000_0000)       
        led <= ~counter1[23:18];
    else if (counter == 32'd1_2500_0000)       
        led <= ~counter1[17:12];
    else if (counter == 32'd1_5000_0000)       
        led <= ~counter1[11:6];
    else if (counter == 32'd1_7500_0000)       
        led <= ~counter1[5:0];
    else if (counter == 32'd2_0000_0000)       
        led <= 6'b000000;
    else if (counter == 32'd2_2500_0000)       
        led <= 6'b111111;
    else if (counter == 32'd2_5000_0000)       
        led <= 6'b000000;
    else
        led <= led;
end
endmodule